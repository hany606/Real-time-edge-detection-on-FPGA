//This implementation of Dual port RAM
//Which has the ability to write and read simultanuosly in different clocks
//This Buffer has two inside ports Buffer A(150x150x8) and B(150x150x1)
module Buffer(
	input [7:0]d_in_a,			// Port A input data
	input [14:0] r_addr_a,		// Port A address for reading
	input [14:0] w_addr_a,		//	Port A address for writing
	input d_in_b,					// Port B input data
	input [14:0] r_addr_b,		//	Port B address for reading
	input [14:0] w_addr_b,		// Port B address for writing
	input w_clk,					//	Write clock (25MHz)
	input r_clk,					//	Read clock  (50MHz)
	input w_en_a,					//	Port A write flag enable
	input w_en_b,					// Port B write flag enable
	output reg [7:0] d_out_a,	// Port A data out (8-bits)
	output reg err_w_a	,		// Port A error in writing
	output reg d_out_b,			// Port A data out (1-bit)
	output reg err_w_b			// Port B error in writing
);

	reg [7:0] data_a[22499:0]; //Registers array (150x150x8) 
	reg data_b[22499:0]; 		//Registers array (150x150x1)
	
	
	//This the initial data for the grayscale static image
	//This was generated by python code to test the algorithm
	initial
	begin
		data_a[0]<=8'd254;
		data_a[1]<=8'd252;
		data_a[2]<=8'd254;
		data_a[3]<=8'd254;
		data_a[4]<=8'd255;
		data_a[5]<=8'd253;
		data_a[6]<=8'd254;
		data_a[7]<=8'd255;
		data_a[8]<=8'd254;
		data_a[9]<=8'd255;
		data_a[10]<=8'd255;
		data_a[11]<=8'd254;
		data_a[12]<=8'd255;
		data_a[13]<=8'd255;
		data_a[14]<=8'd254;
		data_a[15]<=8'd254;
		data_a[16]<=8'd255;
		data_a[17]<=8'd255;
		data_a[18]<=8'd255;
		data_a[19]<=8'd255;
		data_a[20]<=8'd255;
		data_a[21]<=8'd255;
		data_a[22]<=8'd255;
		data_a[23]<=8'd255;
		data_a[24]<=8'd254;
		data_a[25]<=8'd255;
		data_a[26]<=8'd255;
		data_a[27]<=8'd255;
		data_a[28]<=8'd255;
		data_a[29]<=8'd254;
		data_a[30]<=8'd254;
		data_a[31]<=8'd254;
		data_a[32]<=8'd255;
		data_a[33]<=8'd255;
		data_a[34]<=8'd254;
		data_a[35]<=8'd254;
		data_a[36]<=8'd255;
		data_a[37]<=8'd255;
		data_a[38]<=8'd255;
		data_a[39]<=8'd255;
		data_a[40]<=8'd255;
		data_a[41]<=8'd253;
		data_a[42]<=8'd254;
		data_a[43]<=8'd255;
		data_a[44]<=8'd253;
		data_a[45]<=8'd255;
		data_a[46]<=8'd255;
		data_a[47]<=8'd253;
		data_a[48]<=8'd255;
		data_a[49]<=8'd255;
		data_a[50]<=8'd255;
		data_a[51]<=8'd255;
		data_a[52]<=8'd255;
		data_a[53]<=8'd255;
		data_a[54]<=8'd254;
		data_a[55]<=8'd254;
		data_a[56]<=8'd255;
		data_a[57]<=8'd255;
		data_a[58]<=8'd255;
		data_a[59]<=8'd255;
		data_a[60]<=8'd255;
		data_a[61]<=8'd255;
		data_a[62]<=8'd255;
		data_a[63]<=8'd255;
		data_a[64]<=8'd254;
		data_a[65]<=8'd254;
		data_a[66]<=8'd254;
		data_a[67]<=8'd254;
		data_a[68]<=8'd254;
		data_a[69]<=8'd255;
		data_a[70]<=8'd255;
		data_a[71]<=8'd254;
		data_a[72]<=8'd254;
		data_a[73]<=8'd254;
		data_a[74]<=8'd254;
		data_a[75]<=8'd255;
		data_a[76]<=8'd255;
		data_a[77]<=8'd255;
		data_a[78]<=8'd254;
		data_a[79]<=8'd254;
		data_a[80]<=8'd254;
		data_a[81]<=8'd254;
		data_a[82]<=8'd253;
		data_a[83]<=8'd254;
		data_a[84]<=8'd254;
		data_a[85]<=8'd255;
		data_a[86]<=8'd254;
		data_a[87]<=8'd255;
		data_a[88]<=8'd255;
		data_a[89]<=8'd255;
		data_a[90]<=8'd254;
		data_a[91]<=8'd254;
		data_a[92]<=8'd254;
		data_a[93]<=8'd254;
		data_a[94]<=8'd254;
		data_a[95]<=8'd254;
		data_a[96]<=8'd254;
		data_a[97]<=8'd254;
		data_a[98]<=8'd252;
		data_a[99]<=8'd254;
		data_a[100]<=8'd254;
		data_a[101]<=8'd252;
		data_a[102]<=8'd255;
		data_a[103]<=8'd255;
		data_a[104]<=8'd255;
		data_a[105]<=8'd254;
		data_a[106]<=8'd255;
		data_a[107]<=8'd255;
		data_a[108]<=8'd253;
		data_a[109]<=8'd253;
		data_a[110]<=8'd255;
		data_a[111]<=8'd255;
		data_a[112]<=8'd255;
		data_a[113]<=8'd253;
		data_a[114]<=8'd255;
		data_a[115]<=8'd255;
		data_a[116]<=8'd255;
		data_a[117]<=8'd255;
		data_a[118]<=8'd254;
		data_a[119]<=8'd254;
		data_a[120]<=8'd254;
		data_a[121]<=8'd254;
		data_a[122]<=8'd254;
		data_a[123]<=8'd254;
		data_a[124]<=8'd254;
		data_a[125]<=8'd253;
		data_a[126]<=8'd254;
		data_a[127]<=8'd253;
		data_a[128]<=8'd254;
		data_a[129]<=8'd254;
		data_a[130]<=8'd254;
		data_a[131]<=8'd254;
		data_a[132]<=8'd254;
		data_a[133]<=8'd254;
		data_a[134]<=8'd254;
		data_a[135]<=8'd254;
		data_a[136]<=8'd254;
		data_a[137]<=8'd254;
		data_a[138]<=8'd254;
		data_a[139]<=8'd254;
		data_a[140]<=8'd254;
		data_a[141]<=8'd254;
		data_a[142]<=8'd254;
		data_a[143]<=8'd254;
		data_a[144]<=8'd254;
		data_a[145]<=8'd254;
		data_a[146]<=8'd254;
		data_a[147]<=8'd254;
		data_a[148]<=8'd254;
		data_a[149]<=8'd254;
		data_a[150]<=8'd252;
		data_a[151]<=8'd228;
		data_a[152]<=8'd227;
		data_a[153]<=8'd223;
		data_a[154]<=8'd220;
		data_a[155]<=8'd225;
		data_a[156]<=8'd225;
		data_a[157]<=8'd209;
		data_a[158]<=8'd216;
		data_a[159]<=8'd219;
		data_a[160]<=8'd221;
		data_a[161]<=8'd222;
		data_a[162]<=8'd223;
		data_a[163]<=8'd223;
		data_a[164]<=8'd221;
		data_a[165]<=8'd219;
		data_a[166]<=8'd218;
		data_a[167]<=8'd218;
		data_a[168]<=8'd218;
		data_a[169]<=8'd219;
		data_a[170]<=8'd219;
		data_a[171]<=8'd219;
		data_a[172]<=8'd220;
		data_a[173]<=8'd220;
		data_a[174]<=8'd219;
		data_a[175]<=8'd219;
		data_a[176]<=8'd220;
		data_a[177]<=8'd220;
		data_a[178]<=8'd219;
		data_a[179]<=8'd219;
		data_a[180]<=8'd218;
		data_a[181]<=8'd218;
		data_a[182]<=8'd218;
		data_a[183]<=8'd218;
		data_a[184]<=8'd218;
		data_a[185]<=8'd218;
		data_a[186]<=8'd218;
		data_a[187]<=8'd219;
		data_a[188]<=8'd219;
		data_a[189]<=8'd219;
		data_a[190]<=8'd220;
		data_a[191]<=8'd224;
		data_a[192]<=8'd219;
		data_a[193]<=8'd220;
		data_a[194]<=8'd221;
		data_a[195]<=8'd217;
		data_a[196]<=8'd219;
		data_a[197]<=8'd250;
		data_a[198]<=8'd253;
		data_a[199]<=8'd254;
		data_a[200]<=8'd254;
		data_a[201]<=8'd253;
		data_a[202]<=8'd254;
		data_a[203]<=8'd255;
		data_a[204]<=8'd255;
		data_a[205]<=8'd255;
		data_a[206]<=8'd255;
		data_a[207]<=8'd255;
		data_a[208]<=8'd255;
		data_a[209]<=8'd255;
		data_a[210]<=8'd255;
		data_a[211]<=8'd255;
		data_a[212]<=8'd255;
		data_a[213]<=8'd255;
		data_a[214]<=8'd254;
		data_a[215]<=8'd254;
		data_a[216]<=8'd254;
		data_a[217]<=8'd255;
		data_a[218]<=8'd255;
		data_a[219]<=8'd255;
		data_a[220]<=8'd255;
		data_a[221]<=8'd254;
		data_a[222]<=8'd254;
		data_a[223]<=8'd248;
		data_a[224]<=8'd230;
		data_a[225]<=8'd229;
		data_a[226]<=8'd216;
		data_a[227]<=8'd224;
		data_a[228]<=8'd223;
		data_a[229]<=8'd223;
		data_a[230]<=8'd217;
		data_a[231]<=8'd220;
		data_a[232]<=8'd223;
		data_a[233]<=8'd220;
		data_a[234]<=8'd214;
		data_a[235]<=8'd211;
		data_a[236]<=8'd213;
		data_a[237]<=8'd218;
		data_a[238]<=8'd219;
		data_a[239]<=8'd218;
		data_a[240]<=8'd217;
		data_a[241]<=8'd217;
		data_a[242]<=8'd218;
		data_a[243]<=8'd219;
		data_a[244]<=8'd218;
		data_a[245]<=8'd217;
		data_a[246]<=8'd215;
		data_a[247]<=8'd215;
		data_a[248]<=8'd217;
		data_a[249]<=8'd214;
		data_a[250]<=8'd206;
		data_a[251]<=8'd220;
		data_a[252]<=8'd218;
		data_a[253]<=8'd217;
		data_a[254]<=8'd219;
		data_a[255]<=8'd211;
		data_a[256]<=8'd219;
		data_a[257]<=8'd213;
		data_a[258]<=8'd219;
		data_a[259]<=8'd226;
		data_a[260]<=8'd219;
		data_a[261]<=8'd210;
		data_a[262]<=8'd221;
		data_a[263]<=8'd223;
		data_a[264]<=8'd222;
		data_a[265]<=8'd222;
		data_a[266]<=8'd225;
		data_a[267]<=8'd223;
		data_a[268]<=8'd222;
		data_a[269]<=8'd225;
		data_a[270]<=8'd225;
		data_a[271]<=8'd226;
		data_a[272]<=8'd226;
		data_a[273]<=8'd225;
		data_a[274]<=8'd227;
		data_a[275]<=8'd224;
		data_a[276]<=8'd228;
		data_a[277]<=8'd227;
		data_a[278]<=8'd228;
		data_a[279]<=8'd228;
		data_a[280]<=8'd228;
		data_a[281]<=8'd228;
		data_a[282]<=8'd228;
		data_a[283]<=8'd228;
		data_a[284]<=8'd228;
		data_a[285]<=8'd228;
		data_a[286]<=8'd232;
		data_a[287]<=8'd233;
		data_a[288]<=8'd233;
		data_a[289]<=8'd234;
		data_a[290]<=8'd234;
		data_a[291]<=8'd235;
		data_a[292]<=8'd237;
		data_a[293]<=8'd238;
		data_a[294]<=8'd236;
		data_a[295]<=8'd236;
		data_a[296]<=8'd236;
		data_a[297]<=8'd236;
		data_a[298]<=8'd235;
		data_a[299]<=8'd234;
		data_a[300]<=8'd254;
		data_a[301]<=8'd225;
		data_a[302]<=8'd225;
		data_a[303]<=8'd228;
		data_a[304]<=8'd221;
		data_a[305]<=8'd209;
		data_a[306]<=8'd209;
		data_a[307]<=8'd222;
		data_a[308]<=8'd220;
		data_a[309]<=8'd222;
		data_a[310]<=8'd222;
		data_a[311]<=8'd221;
		data_a[312]<=8'd220;
		data_a[313]<=8'd220;
		data_a[314]<=8'd220;
		data_a[315]<=8'd220;
		data_a[316]<=8'd217;
		data_a[317]<=8'd218;
		data_a[318]<=8'd218;
		data_a[319]<=8'd218;
		data_a[320]<=8'd219;
		data_a[321]<=8'd219;
		data_a[322]<=8'd220;
		data_a[323]<=8'd220;
		data_a[324]<=8'd219;
		data_a[325]<=8'd219;
		data_a[326]<=8'd218;
		data_a[327]<=8'd218;
		data_a[328]<=8'd218;
		data_a[329]<=8'd218;
		data_a[330]<=8'd218;
		data_a[331]<=8'd218;
		data_a[332]<=8'd218;
		data_a[333]<=8'd218;
		data_a[334]<=8'd218;
		data_a[335]<=8'd217;
		data_a[336]<=8'd218;
		data_a[337]<=8'd218;
		data_a[338]<=8'd218;
		data_a[339]<=8'd219;
		data_a[340]<=8'd220;
		data_a[341]<=8'd221;
		data_a[342]<=8'd223;
		data_a[343]<=8'd221;
		data_a[344]<=8'd219;
		data_a[345]<=8'd231;
		data_a[346]<=8'd224;
		data_a[347]<=8'd209;
		data_a[348]<=8'd255;
		data_a[349]<=8'd255;
		data_a[350]<=8'd255;
		data_a[351]<=8'd255;
		data_a[352]<=8'd255;
		data_a[353]<=8'd254;
		data_a[354]<=8'd254;
		data_a[355]<=8'd255;
		data_a[356]<=8'd255;
		data_a[357]<=8'd255;
		data_a[358]<=8'd255;
		data_a[359]<=8'd255;
		data_a[360]<=8'd255;
		data_a[361]<=8'd255;
		data_a[362]<=8'd255;
		data_a[363]<=8'd255;
		data_a[364]<=8'd254;
		data_a[365]<=8'd254;
		data_a[366]<=8'd254;
		data_a[367]<=8'd255;
		data_a[368]<=8'd255;
		data_a[369]<=8'd255;
		data_a[370]<=8'd255;
		data_a[371]<=8'd254;
		data_a[372]<=8'd252;
		data_a[373]<=8'd254;
		data_a[374]<=8'd221;
		data_a[375]<=8'd228;
		data_a[376]<=8'd225;
		data_a[377]<=8'd222;
		data_a[378]<=8'd221;
		data_a[379]<=8'd221;
		data_a[380]<=8'd222;
		data_a[381]<=8'd217;
		data_a[382]<=8'd211;
		data_a[383]<=8'd210;
		data_a[384]<=8'd214;
		data_a[385]<=8'd219;
		data_a[386]<=8'd218;
		data_a[387]<=8'd216;
		data_a[388]<=8'd218;
		data_a[389]<=8'd216;
		data_a[390]<=8'd215;
		data_a[391]<=8'd216;
		data_a[392]<=8'd217;
		data_a[393]<=8'd218;
		data_a[394]<=8'd217;
		data_a[395]<=8'd217;
		data_a[396]<=8'd216;
		data_a[397]<=8'd211;
		data_a[398]<=8'd218;
		data_a[399]<=8'd216;
		data_a[400]<=8'd207;
		data_a[401]<=8'd217;
		data_a[402]<=8'd219;
		data_a[403]<=8'd218;
		data_a[404]<=8'd215;
		data_a[405]<=8'd226;
		data_a[406]<=8'd220;
		data_a[407]<=8'd207;
		data_a[408]<=8'd213;
		data_a[409]<=8'd215;
		data_a[410]<=8'd216;
		data_a[411]<=8'd225;
		data_a[412]<=8'd218;
		data_a[413]<=8'd223;
		data_a[414]<=8'd221;
		data_a[415]<=8'd220;
		data_a[416]<=8'd226;
		data_a[417]<=8'd224;
		data_a[418]<=8'd221;
		data_a[419]<=8'd227;
		data_a[420]<=8'd225;
		data_a[421]<=8'd226;
		data_a[422]<=8'd226;
		data_a[423]<=8'd225;
		data_a[424]<=8'd227;
		data_a[425]<=8'd224;
		data_a[426]<=8'd229;
		data_a[427]<=8'd228;
		data_a[428]<=8'd229;
		data_a[429]<=8'd229;
		data_a[430]<=8'd229;
		data_a[431]<=8'd230;
		data_a[432]<=8'd230;
		data_a[433]<=8'd230;
		data_a[434]<=8'd230;
		data_a[435]<=8'd230;
		data_a[436]<=8'd230;
		data_a[437]<=8'd231;
		data_a[438]<=8'd232;
		data_a[439]<=8'd233;
		data_a[440]<=8'd233;
		data_a[441]<=8'd235;
		data_a[442]<=8'd237;
		data_a[443]<=8'd239;
		data_a[444]<=8'd238;
		data_a[445]<=8'd239;
		data_a[446]<=8'd240;
		data_a[447]<=8'd239;
		data_a[448]<=8'd237;
		data_a[449]<=8'd235;
		data_a[450]<=8'd251;
		data_a[451]<=8'd230;
		data_a[452]<=8'd228;
		data_a[453]<=8'd216;
		data_a[454]<=8'd216;
		data_a[455]<=8'd225;
		data_a[456]<=8'd222;
		data_a[457]<=8'd220;
		data_a[458]<=8'd224;
		data_a[459]<=8'd224;
		data_a[460]<=8'd223;
		data_a[461]<=8'd221;
		data_a[462]<=8'd219;
		data_a[463]<=8'd219;
		data_a[464]<=8'd220;
		data_a[465]<=8'd221;
		data_a[466]<=8'd219;
		data_a[467]<=8'd219;
		data_a[468]<=8'd220;
		data_a[469]<=8'd220;
		data_a[470]<=8'd220;
		data_a[471]<=8'd220;
		data_a[472]<=8'd220;
		data_a[473]<=8'd220;
		data_a[474]<=8'd221;
		data_a[475]<=8'd220;
		data_a[476]<=8'd218;
		data_a[477]<=8'd218;
		data_a[478]<=8'd219;
		data_a[479]<=8'd219;
		data_a[480]<=8'd219;
		data_a[481]<=8'd219;
		data_a[482]<=8'd219;
		data_a[483]<=8'd219;
		data_a[484]<=8'd218;
		data_a[485]<=8'd218;
		data_a[486]<=8'd218;
		data_a[487]<=8'd219;
		data_a[488]<=8'd219;
		data_a[489]<=8'd219;
		data_a[490]<=8'd217;
		data_a[491]<=8'd216;
		data_a[492]<=8'd218;
		data_a[493]<=8'd222;
		data_a[494]<=8'd223;
		data_a[495]<=8'd221;
		data_a[496]<=8'd224;
		data_a[497]<=8'd239;
		data_a[498]<=8'd244;
		data_a[499]<=8'd249;
		data_a[500]<=8'd253;
		data_a[501]<=8'd255;
		data_a[502]<=8'd254;
		data_a[503]<=8'd254;
		data_a[504]<=8'd254;
		data_a[505]<=8'd254;
		data_a[506]<=8'd255;
		data_a[507]<=8'd255;
		data_a[508]<=8'd255;
		data_a[509]<=8'd255;
		data_a[510]<=8'd255;
		data_a[511]<=8'd255;
		data_a[512]<=8'd255;
		data_a[513]<=8'd255;
		data_a[514]<=8'd254;
		data_a[515]<=8'd254;
		data_a[516]<=8'd254;
		data_a[517]<=8'd255;
		data_a[518]<=8'd255;
		data_a[519]<=8'd255;
		data_a[520]<=8'd255;
		data_a[521]<=8'd254;
		data_a[522]<=8'd254;
		data_a[523]<=8'd251;
		data_a[524]<=8'd242;
		data_a[525]<=8'd230;
		data_a[526]<=8'd223;
		data_a[527]<=8'd221;
		data_a[528]<=8'd227;
		data_a[529]<=8'd221;
		data_a[530]<=8'd213;
		data_a[531]<=8'd215;
		data_a[532]<=8'd217;
		data_a[533]<=8'd220;
		data_a[534]<=8'd223;
		data_a[535]<=8'd224;
		data_a[536]<=8'd220;
		data_a[537]<=8'd215;
		data_a[538]<=8'd218;
		data_a[539]<=8'd217;
		data_a[540]<=8'd216;
		data_a[541]<=8'd217;
		data_a[542]<=8'd218;
		data_a[543]<=8'd218;
		data_a[544]<=8'd218;
		data_a[545]<=8'd218;
		data_a[546]<=8'd215;
		data_a[547]<=8'd213;
		data_a[548]<=8'd218;
		data_a[549]<=8'd217;
		data_a[550]<=8'd219;
		data_a[551]<=8'd207;
		data_a[552]<=8'd217;
		data_a[553]<=8'd210;
		data_a[554]<=8'd219;
		data_a[555]<=8'd193;
		data_a[556]<=8'd190;
		data_a[557]<=8'd151;
		data_a[558]<=8'd232;
		data_a[559]<=8'd225;
		data_a[560]<=8'd216;
		data_a[561]<=8'd218;
		data_a[562]<=8'd218;
		data_a[563]<=8'd222;
		data_a[564]<=8'd220;
		data_a[565]<=8'd220;
		data_a[566]<=8'd225;
		data_a[567]<=8'd223;
		data_a[568]<=8'd221;
		data_a[569]<=8'd226;
		data_a[570]<=8'd223;
		data_a[571]<=8'd224;
		data_a[572]<=8'd224;
		data_a[573]<=8'd223;
		data_a[574]<=8'd226;
		data_a[575]<=8'd223;
		data_a[576]<=8'd227;
		data_a[577]<=8'd226;
		data_a[578]<=8'd227;
		data_a[579]<=8'd227;
		data_a[580]<=8'd228;
		data_a[581]<=8'd229;
		data_a[582]<=8'd229;
		data_a[583]<=8'd229;
		data_a[584]<=8'd230;
		data_a[585]<=8'd230;
		data_a[586]<=8'd234;
		data_a[587]<=8'd235;
		data_a[588]<=8'd237;
		data_a[589]<=8'd237;
		data_a[590]<=8'd236;
		data_a[591]<=8'd237;
		data_a[592]<=8'd239;
		data_a[593]<=8'd241;
		data_a[594]<=8'd238;
		data_a[595]<=8'd239;
		data_a[596]<=8'd239;
		data_a[597]<=8'd239;
		data_a[598]<=8'd238;
		data_a[599]<=8'd237;
		data_a[600]<=8'd255;
		data_a[601]<=8'd218;
		data_a[602]<=8'd221;
		data_a[603]<=8'd224;
		data_a[604]<=8'd221;
		data_a[605]<=8'd226;
		data_a[606]<=8'd226;
		data_a[607]<=8'd221;
		data_a[608]<=8'd220;
		data_a[609]<=8'd222;
		data_a[610]<=8'd223;
		data_a[611]<=8'd223;
		data_a[612]<=8'd222;
		data_a[613]<=8'd220;
		data_a[614]<=8'd219;
		data_a[615]<=8'd219;
		data_a[616]<=8'd220;
		data_a[617]<=8'd220;
		data_a[618]<=8'd220;
		data_a[619]<=8'd220;
		data_a[620]<=8'd219;
		data_a[621]<=8'd219;
		data_a[622]<=8'd219;
		data_a[623]<=8'd218;
		data_a[624]<=8'd220;
		data_a[625]<=8'd219;
		data_a[626]<=8'd217;
		data_a[627]<=8'd217;
		data_a[628]<=8'd218;
		data_a[629]<=8'd218;
		data_a[630]<=8'd218;
		data_a[631]<=8'd218;
		data_a[632]<=8'd218;
		data_a[633]<=8'd218;
		data_a[634]<=8'd218;
		data_a[635]<=8'd218;
		data_a[636]<=8'd218;
		data_a[637]<=8'd218;
		data_a[638]<=8'd218;
		data_a[639]<=8'd218;
		data_a[640]<=8'd220;
		data_a[641]<=8'd223;
		data_a[642]<=8'd224;
		data_a[643]<=8'd219;
		data_a[644]<=8'd221;
		data_a[645]<=8'd227;
		data_a[646]<=8'd228;
		data_a[647]<=8'd227;
		data_a[648]<=8'd228;
		data_a[649]<=8'd243;
		data_a[650]<=8'd254;
		data_a[651]<=8'd253;
		data_a[652]<=8'd253;
		data_a[653]<=8'd255;
		data_a[654]<=8'd255;
		data_a[655]<=8'd253;
		data_a[656]<=8'd255;
		data_a[657]<=8'd255;
		data_a[658]<=8'd255;
		data_a[659]<=8'd255;
		data_a[660]<=8'd255;
		data_a[661]<=8'd255;
		data_a[662]<=8'd255;
		data_a[663]<=8'd255;
		data_a[664]<=8'd254;
		data_a[665]<=8'd254;
		data_a[666]<=8'd255;
		data_a[667]<=8'd255;
		data_a[668]<=8'd255;
		data_a[669]<=8'd255;
		data_a[670]<=8'd255;
		data_a[671]<=8'd255;
		data_a[672]<=8'd254;
		data_a[673]<=8'd255;
		data_a[674]<=8'd255;
		data_a[675]<=8'd214;
		data_a[676]<=8'd219;
		data_a[677]<=8'd228;
		data_a[678]<=8'd211;
		data_a[679]<=8'd214;
		data_a[680]<=8'd218;
		data_a[681]<=8'd221;
		data_a[682]<=8'd222;
		data_a[683]<=8'd219;
		data_a[684]<=8'd216;
		data_a[685]<=8'd216;
		data_a[686]<=8'd218;
		data_a[687]<=8'd219;
		data_a[688]<=8'd218;
		data_a[689]<=8'd216;
		data_a[690]<=8'd215;
		data_a[691]<=8'd216;
		data_a[692]<=8'd217;
		data_a[693]<=8'd216;
		data_a[694]<=8'd216;
		data_a[695]<=8'd216;
		data_a[696]<=8'd212;
		data_a[697]<=8'd218;
		data_a[698]<=8'd218;
		data_a[699]<=8'd213;
		data_a[700]<=8'd220;
		data_a[701]<=8'd208;
		data_a[702]<=8'd212;
		data_a[703]<=8'd206;
		data_a[704]<=8'd209;
		data_a[705]<=8'd219;
		data_a[706]<=8'd215;
		data_a[707]<=8'd196;
		data_a[708]<=8'd159;
		data_a[709]<=8'd191;
		data_a[710]<=8'd220;
		data_a[711]<=8'd221;
		data_a[712]<=8'd221;
		data_a[713]<=8'd220;
		data_a[714]<=8'd221;
		data_a[715]<=8'd223;
		data_a[716]<=8'd223;
		data_a[717]<=8'd223;
		data_a[718]<=8'd223;
		data_a[719]<=8'd223;
		data_a[720]<=8'd223;
		data_a[721]<=8'd224;
		data_a[722]<=8'd225;
		data_a[723]<=8'd225;
		data_a[724]<=8'd227;
		data_a[725]<=8'd223;
		data_a[726]<=8'd227;
		data_a[727]<=8'd225;
		data_a[728]<=8'd227;
		data_a[729]<=8'd228;
		data_a[730]<=8'd229;
		data_a[731]<=8'd230;
		data_a[732]<=8'd230;
		data_a[733]<=8'd231;
		data_a[734]<=8'd232;
		data_a[735]<=8'd232;
		data_a[736]<=8'd233;
		data_a[737]<=8'd235;
		data_a[738]<=8'd237;
		data_a[739]<=8'd237;
		data_a[740]<=8'd236;
		data_a[741]<=8'd236;
		data_a[742]<=8'd238;
		data_a[743]<=8'd240;
		data_a[744]<=8'd241;
		data_a[745]<=8'd241;
		data_a[746]<=8'd240;
		data_a[747]<=8'd240;
		data_a[748]<=8'd241;
		data_a[749]<=8'd241;
		data_a[750]<=8'd254;
		data_a[751]<=8'd223;
		data_a[752]<=8'd226;
		data_a[753]<=8'd228;
		data_a[754]<=8'd224;
		data_a[755]<=8'd221;
		data_a[756]<=8'd222;
		data_a[757]<=8'd225;
		data_a[758]<=8'd222;
		data_a[759]<=8'd222;
		data_a[760]<=8'd222;
		data_a[761]<=8'd221;
		data_a[762]<=8'd220;
		data_a[763]<=8'd218;
		data_a[764]<=8'd218;
		data_a[765]<=8'd219;
		data_a[766]<=8'd220;
		data_a[767]<=8'd220;
		data_a[768]<=8'd220;
		data_a[769]<=8'd220;
		data_a[770]<=8'd219;
		data_a[771]<=8'd219;
		data_a[772]<=8'd218;
		data_a[773]<=8'd217;
		data_a[774]<=8'd219;
		data_a[775]<=8'd218;
		data_a[776]<=8'd218;
		data_a[777]<=8'd218;
		data_a[778]<=8'd218;
		data_a[779]<=8'd218;
		data_a[780]<=8'd218;
		data_a[781]<=8'd217;
		data_a[782]<=8'd218;
		data_a[783]<=8'd218;
		data_a[784]<=8'd218;
		data_a[785]<=8'd217;
		data_a[786]<=8'd217;
		data_a[787]<=8'd218;
		data_a[788]<=8'd218;
		data_a[789]<=8'd218;
		data_a[790]<=8'd217;
		data_a[791]<=8'd221;
		data_a[792]<=8'd219;
		data_a[793]<=8'd213;
		data_a[794]<=8'd223;
		data_a[795]<=8'd224;
		data_a[796]<=8'd224;
		data_a[797]<=8'd234;
		data_a[798]<=8'd227;
		data_a[799]<=8'd235;
		data_a[800]<=8'd247;
		data_a[801]<=8'd255;
		data_a[802]<=8'd255;
		data_a[803]<=8'd255;
		data_a[804]<=8'd254;
		data_a[805]<=8'd255;
		data_a[806]<=8'd255;
		data_a[807]<=8'd255;
		data_a[808]<=8'd255;
		data_a[809]<=8'd255;
		data_a[810]<=8'd255;
		data_a[811]<=8'd255;
		data_a[812]<=8'd255;
		data_a[813]<=8'd255;
		data_a[814]<=8'd254;
		data_a[815]<=8'd255;
		data_a[816]<=8'd255;
		data_a[817]<=8'd255;
		data_a[818]<=8'd255;
		data_a[819]<=8'd255;
		data_a[820]<=8'd255;
		data_a[821]<=8'd255;
		data_a[822]<=8'd252;
		data_a[823]<=8'd255;
		data_a[824]<=8'd251;
		data_a[825]<=8'd231;
		data_a[826]<=8'd216;
		data_a[827]<=8'd217;
		data_a[828]<=8'd219;
		data_a[829]<=8'd222;
		data_a[830]<=8'd219;
		data_a[831]<=8'd219;
		data_a[832]<=8'd220;
		data_a[833]<=8'd221;
		data_a[834]<=8'd221;
		data_a[835]<=8'd220;
		data_a[836]<=8'd216;
		data_a[837]<=8'd212;
		data_a[838]<=8'd219;
		data_a[839]<=8'd217;
		data_a[840]<=8'd215;
		data_a[841]<=8'd216;
		data_a[842]<=8'd216;
		data_a[843]<=8'd214;
		data_a[844]<=8'd213;
		data_a[845]<=8'd214;
		data_a[846]<=8'd215;
		data_a[847]<=8'd216;
		data_a[848]<=8'd215;
		data_a[849]<=8'd214;
		data_a[850]<=8'd218;
		data_a[851]<=8'd218;
		data_a[852]<=8'd208;
		data_a[853]<=8'd219;
		data_a[854]<=8'd213;
		data_a[855]<=8'd211;
		data_a[856]<=8'd220;
		data_a[857]<=8'd215;
		data_a[858]<=8'd211;
		data_a[859]<=8'd180;
		data_a[860]<=8'd179;
		data_a[861]<=8'd223;
		data_a[862]<=8'd220;
		data_a[863]<=8'd218;
		data_a[864]<=8'd221;
		data_a[865]<=8'd224;
		data_a[866]<=8'd222;
		data_a[867]<=8'd222;
		data_a[868]<=8'd223;
		data_a[869]<=8'd221;
		data_a[870]<=8'd222;
		data_a[871]<=8'd224;
		data_a[872]<=8'd225;
		data_a[873]<=8'd224;
		data_a[874]<=8'd226;
		data_a[875]<=8'd222;
		data_a[876]<=8'd226;
		data_a[877]<=8'd225;
		data_a[878]<=8'd227;
		data_a[879]<=8'd228;
		data_a[880]<=8'd230;
		data_a[881]<=8'd230;
		data_a[882]<=8'd231;
		data_a[883]<=8'd232;
		data_a[884]<=8'd233;
		data_a[885]<=8'd234;
		data_a[886]<=8'd235;
		data_a[887]<=8'd236;
		data_a[888]<=8'd239;
		data_a[889]<=8'd240;
		data_a[890]<=8'd240;
		data_a[891]<=8'd240;
		data_a[892]<=8'd242;
		data_a[893]<=8'd243;
		data_a[894]<=8'd242;
		data_a[895]<=8'd241;
		data_a[896]<=8'd241;
		data_a[897]<=8'd241;
		data_a[898]<=8'd243;
		data_a[899]<=8'd244;
		data_a[900]<=8'd254;
		data_a[901]<=8'd234;
		data_a[902]<=8'd228;
		data_a[903]<=8'd227;
		data_a[904]<=8'd232;
		data_a[905]<=8'd226;
		data_a[906]<=8'd222;
		data_a[907]<=8'd225;
		data_a[908]<=8'd225;
		data_a[909]<=8'd223;
		data_a[910]<=8'd220;
		data_a[911]<=8'd219;
		data_a[912]<=8'd217;
		data_a[913]<=8'd217;
		data_a[914]<=8'd218;
		data_a[915]<=8'd220;
		data_a[916]<=8'd219;
		data_a[917]<=8'd220;
		data_a[918]<=8'd220;
		data_a[919]<=8'd220;
		data_a[920]<=8'd220;
		data_a[921]<=8'd219;
		data_a[922]<=8'd218;
		data_a[923]<=8'd218;
		data_a[924]<=8'd218;
		data_a[925]<=8'd219;
		data_a[926]<=8'd219;
		data_a[927]<=8'd219;
		data_a[928]<=8'd219;
		data_a[929]<=8'd218;
		data_a[930]<=8'd218;
		data_a[931]<=8'd218;
		data_a[932]<=8'd218;
		data_a[933]<=8'd218;
		data_a[934]<=8'd218;
		data_a[935]<=8'd218;
		data_a[936]<=8'd218;
		data_a[937]<=8'd218;
		data_a[938]<=8'd218;
		data_a[939]<=8'd218;
		data_a[940]<=8'd222;
		data_a[941]<=8'd211;
		data_a[942]<=8'd220;
		data_a[943]<=8'd223;
		data_a[944]<=8'd222;
		data_a[945]<=8'd222;
		data_a[946]<=8'd227;
		data_a[947]<=8'd224;
		data_a[948]<=8'd224;
		data_a[949]<=8'd224;
		data_a[950]<=8'd234;
		data_a[951]<=8'd251;
		data_a[952]<=8'd255;
		data_a[953]<=8'd253;
		data_a[954]<=8'd252;
		data_a[955]<=8'd255;
		data_a[956]<=8'd255;
		data_a[957]<=8'd255;
		data_a[958]<=8'd255;
		data_a[959]<=8'd255;
		data_a[960]<=8'd255;
		data_a[961]<=8'd255;
		data_a[962]<=8'd255;
		data_a[963]<=8'd255;
		data_a[964]<=8'd254;
		data_a[965]<=8'd255;
		data_a[966]<=8'd255;
		data_a[967]<=8'd255;
		data_a[968]<=8'd255;
		data_a[969]<=8'd253;
		data_a[970]<=8'd252;
		data_a[971]<=8'd251;
		data_a[972]<=8'd248;
		data_a[973]<=8'd252;
		data_a[974]<=8'd215;
		data_a[975]<=8'd222;
		data_a[976]<=8'd225;
		data_a[977]<=8'd218;
		data_a[978]<=8'd219;
		data_a[979]<=8'd220;
		data_a[980]<=8'd220;
		data_a[981]<=8'd219;
		data_a[982]<=8'd219;
		data_a[983]<=8'd218;
		data_a[984]<=8'd217;
		data_a[985]<=8'd217;
		data_a[986]<=8'd219;
		data_a[987]<=8'd221;
		data_a[988]<=8'd218;
		data_a[989]<=8'd216;
		data_a[990]<=8'd215;
		data_a[991]<=8'd216;
		data_a[992]<=8'd215;
		data_a[993]<=8'd214;
		data_a[994]<=8'd213;
		data_a[995]<=8'd214;
		data_a[996]<=8'd214;
		data_a[997]<=8'd212;
		data_a[998]<=8'd211;
		data_a[999]<=8'd216;
		data_a[1000]<=8'd214;
		data_a[1001]<=8'd216;
		data_a[1002]<=8'd208;
		data_a[1003]<=8'd222;
		data_a[1004]<=8'd218;
		data_a[1005]<=8'd221;
		data_a[1006]<=8'd216;
		data_a[1007]<=8'd213;
		data_a[1008]<=8'd204;
		data_a[1009]<=8'd218;
		data_a[1010]<=8'd219;
		data_a[1011]<=8'd184;
		data_a[1012]<=8'd214;
		data_a[1013]<=8'd217;
		data_a[1014]<=8'd220;
		data_a[1015]<=8'd222;
		data_a[1016]<=8'd221;
		data_a[1017]<=8'd220;
		data_a[1018]<=8'd220;
		data_a[1019]<=8'd222;
		data_a[1020]<=8'd220;
		data_a[1021]<=8'd222;
		data_a[1022]<=8'd223;
		data_a[1023]<=8'd222;
		data_a[1024]<=8'd224;
		data_a[1025]<=8'd220;
		data_a[1026]<=8'd225;
		data_a[1027]<=8'd224;
		data_a[1028]<=8'd225;
		data_a[1029]<=8'd227;
		data_a[1030]<=8'd229;
		data_a[1031]<=8'd230;
		data_a[1032]<=8'd230;
		data_a[1033]<=8'd231;
		data_a[1034]<=8'd233;
		data_a[1035]<=8'd234;
		data_a[1036]<=8'd235;
		data_a[1037]<=8'd236;
		data_a[1038]<=8'd237;
		data_a[1039]<=8'd239;
		data_a[1040]<=8'd240;
		data_a[1041]<=8'd242;
		data_a[1042]<=8'd243;
		data_a[1043]<=8'd244;
		data_a[1044]<=8'd247;
		data_a[1045]<=8'd247;
		data_a[1046]<=8'd247;
		data_a[1047]<=8'd248;
		data_a[1048]<=8'd248;
		data_a[1049]<=8'd249;
		data_a[1050]<=8'd254;
		data_a[1051]<=8'd234;
		data_a[1052]<=8'd229;
		data_a[1053]<=8'd228;
		data_a[1054]<=8'd226;
		data_a[1055]<=8'd223;
		data_a[1056]<=8'd225;
		data_a[1057]<=8'd220;
		data_a[1058]<=8'd222;
		data_a[1059]<=8'd220;
		data_a[1060]<=8'd220;
		data_a[1061]<=8'd221;
		data_a[1062]<=8'd220;
		data_a[1063]<=8'd219;
		data_a[1064]<=8'd218;
		data_a[1065]<=8'd219;
		data_a[1066]<=8'd217;
		data_a[1067]<=8'd218;
		data_a[1068]<=8'd218;
		data_a[1069]<=8'd218;
		data_a[1070]<=8'd218;
		data_a[1071]<=8'd218;
		data_a[1072]<=8'd218;
		data_a[1073]<=8'd217;
		data_a[1074]<=8'd217;
		data_a[1075]<=8'd218;
		data_a[1076]<=8'd220;
		data_a[1077]<=8'd220;
		data_a[1078]<=8'd219;
		data_a[1079]<=8'd218;
		data_a[1080]<=8'd217;
		data_a[1081]<=8'd217;
		data_a[1082]<=8'd217;
		data_a[1083]<=8'd217;
		data_a[1084]<=8'd217;
		data_a[1085]<=8'd216;
		data_a[1086]<=8'd216;
		data_a[1087]<=8'd216;
		data_a[1088]<=8'd217;
		data_a[1089]<=8'd217;
		data_a[1090]<=8'd216;
		data_a[1091]<=8'd218;
		data_a[1092]<=8'd222;
		data_a[1093]<=8'd218;
		data_a[1094]<=8'd225;
		data_a[1095]<=8'd218;
		data_a[1096]<=8'd214;
		data_a[1097]<=8'd221;
		data_a[1098]<=8'd231;
		data_a[1099]<=8'd234;
		data_a[1100]<=8'd238;
		data_a[1101]<=8'd245;
		data_a[1102]<=8'd253;
		data_a[1103]<=8'd255;
		data_a[1104]<=8'd255;
		data_a[1105]<=8'd252;
		data_a[1106]<=8'd255;
		data_a[1107]<=8'd255;
		data_a[1108]<=8'd255;
		data_a[1109]<=8'd255;
		data_a[1110]<=8'd255;
		data_a[1111]<=8'd255;
		data_a[1112]<=8'd255;
		data_a[1113]<=8'd255;
		data_a[1114]<=8'd253;
		data_a[1115]<=8'd254;
		data_a[1116]<=8'd255;
		data_a[1117]<=8'd255;
		data_a[1118]<=8'd255;
		data_a[1119]<=8'd252;
		data_a[1120]<=8'd250;
		data_a[1121]<=8'd248;
		data_a[1122]<=8'd213;
		data_a[1123]<=8'd229;
		data_a[1124]<=8'd225;
		data_a[1125]<=8'd225;
		data_a[1126]<=8'd219;
		data_a[1127]<=8'd221;
		data_a[1128]<=8'd217;
		data_a[1129]<=8'd222;
		data_a[1130]<=8'd221;
		data_a[1131]<=8'd219;
		data_a[1132]<=8'd219;
		data_a[1133]<=8'd220;
		data_a[1134]<=8'd219;
		data_a[1135]<=8'd216;
		data_a[1136]<=8'd215;
		data_a[1137]<=8'd216;
		data_a[1138]<=8'd215;
		data_a[1139]<=8'd213;
		data_a[1140]<=8'd213;
		data_a[1141]<=8'd215;
		data_a[1142]<=8'd215;
		data_a[1143]<=8'd214;
		data_a[1144]<=8'd214;
		data_a[1145]<=8'd216;
		data_a[1146]<=8'd212;
		data_a[1147]<=8'd218;
		data_a[1148]<=8'd216;
		data_a[1149]<=8'd215;
		data_a[1150]<=8'd212;
		data_a[1151]<=8'd210;
		data_a[1152]<=8'd214;
		data_a[1153]<=8'd208;
		data_a[1154]<=8'd213;
		data_a[1155]<=8'd215;
		data_a[1156]<=8'd218;
		data_a[1157]<=8'd205;
		data_a[1158]<=8'd209;
		data_a[1159]<=8'd201;
		data_a[1160]<=8'd214;
		data_a[1161]<=8'd204;
		data_a[1162]<=8'd209;
		data_a[1163]<=8'd218;
		data_a[1164]<=8'd220;
		data_a[1165]<=8'd220;
		data_a[1166]<=8'd223;
		data_a[1167]<=8'd219;
		data_a[1168]<=8'd217;
		data_a[1169]<=8'd225;
		data_a[1170]<=8'd220;
		data_a[1171]<=8'd222;
		data_a[1172]<=8'd223;
		data_a[1173]<=8'd222;
		data_a[1174]<=8'd224;
		data_a[1175]<=8'd221;
		data_a[1176]<=8'd226;
		data_a[1177]<=8'd226;
		data_a[1178]<=8'd225;
		data_a[1179]<=8'd227;
		data_a[1180]<=8'd229;
		data_a[1181]<=8'd230;
		data_a[1182]<=8'd231;
		data_a[1183]<=8'd232;
		data_a[1184]<=8'd234;
		data_a[1185]<=8'd235;
		data_a[1186]<=8'd239;
		data_a[1187]<=8'd239;
		data_a[1188]<=8'd240;
		data_a[1189]<=8'd241;
		data_a[1190]<=8'd243;
		data_a[1191]<=8'd245;
		data_a[1192]<=8'd247;
		data_a[1193]<=8'd248;
		data_a[1194]<=8'd251;
		data_a[1195]<=8'd252;
		data_a[1196]<=8'd253;
		data_a[1197]<=8'd254;
		data_a[1198]<=8'd253;
		data_a[1199]<=8'd253;
		data_a[1200]<=8'd254;
		data_a[1201]<=8'd237;
		data_a[1202]<=8'd226;
		data_a[1203]<=8'd228;
		data_a[1204]<=8'd224;
		data_a[1205]<=8'd222;
		data_a[1206]<=8'd222;
		data_a[1207]<=8'd221;
		data_a[1208]<=8'd223;
		data_a[1209]<=8'd223;
		data_a[1210]<=8'd221;
		data_a[1211]<=8'd220;
		data_a[1212]<=8'd219;
		data_a[1213]<=8'd219;
		data_a[1214]<=8'd219;
		data_a[1215]<=8'd219;
		data_a[1216]<=8'd219;
		data_a[1217]<=8'd218;
		data_a[1218]<=8'd217;
		data_a[1219]<=8'd217;
		data_a[1220]<=8'd218;
		data_a[1221]<=8'd218;
		data_a[1222]<=8'd217;
		data_a[1223]<=8'd217;
		data_a[1224]<=8'd219;
		data_a[1225]<=8'd217;
		data_a[1226]<=8'd217;
		data_a[1227]<=8'd219;
		data_a[1228]<=8'd218;
		data_a[1229]<=8'd216;
		data_a[1230]<=8'd216;
		data_a[1231]<=8'd218;
		data_a[1232]<=8'd215;
		data_a[1233]<=8'd217;
		data_a[1234]<=8'd219;
		data_a[1235]<=8'd213;
		data_a[1236]<=8'd215;
		data_a[1237]<=8'd215;
		data_a[1238]<=8'd218;
		data_a[1239]<=8'd214;
		data_a[1240]<=8'd220;
		data_a[1241]<=8'd222;
		data_a[1242]<=8'd218;
		data_a[1243]<=8'd211;
		data_a[1244]<=8'd212;
		data_a[1245]<=8'd221;
		data_a[1246]<=8'd226;
		data_a[1247]<=8'd224;
		data_a[1248]<=8'd229;
		data_a[1249]<=8'd236;
		data_a[1250]<=8'd235;
		data_a[1251]<=8'd237;
		data_a[1252]<=8'd239;
		data_a[1253]<=8'd252;
		data_a[1254]<=8'd254;
		data_a[1255]<=8'd254;
		data_a[1256]<=8'd255;
		data_a[1257]<=8'd255;
		data_a[1258]<=8'd255;
		data_a[1259]<=8'd255;
		data_a[1260]<=8'd255;
		data_a[1261]<=8'd255;
		data_a[1262]<=8'd255;
		data_a[1263]<=8'd255;
		data_a[1264]<=8'd254;
		data_a[1265]<=8'd255;
		data_a[1266]<=8'd255;
		data_a[1267]<=8'd253;
		data_a[1268]<=8'd247;
		data_a[1269]<=8'd240;
		data_a[1270]<=8'd235;
		data_a[1271]<=8'd233;
		data_a[1272]<=8'd228;
		data_a[1273]<=8'd226;
		data_a[1274]<=8'd224;
		data_a[1275]<=8'd221;
		data_a[1276]<=8'd219;
		data_a[1277]<=8'd219;
		data_a[1278]<=8'd220;
		data_a[1279]<=8'd221;
		data_a[1280]<=8'd219;
		data_a[1281]<=8'd217;
		data_a[1282]<=8'd213;
		data_a[1283]<=8'd223;
		data_a[1284]<=8'd211;
		data_a[1285]<=8'd214;
		data_a[1286]<=8'd218;
		data_a[1287]<=8'd218;
		data_a[1288]<=8'd216;
		data_a[1289]<=8'd212;
		data_a[1290]<=8'd220;
		data_a[1291]<=8'd213;
		data_a[1292]<=8'd213;
		data_a[1293]<=8'd217;
		data_a[1294]<=8'd211;
		data_a[1295]<=8'd217;
		data_a[1296]<=8'd212;
		data_a[1297]<=8'd218;
		data_a[1298]<=8'd215;
		data_a[1299]<=8'd214;
		data_a[1300]<=8'd217;
		data_a[1301]<=8'd221;
		data_a[1302]<=8'd220;
		data_a[1303]<=8'd207;
		data_a[1304]<=8'd208;
		data_a[1305]<=8'd218;
		data_a[1306]<=8'd200;
		data_a[1307]<=8'd193;
		data_a[1308]<=8'd179;
		data_a[1309]<=8'd201;
		data_a[1310]<=8'd188;
		data_a[1311]<=8'd211;
		data_a[1312]<=8'd181;
		data_a[1313]<=8'd219;
		data_a[1314]<=8'd227;
		data_a[1315]<=8'd213;
		data_a[1316]<=8'd219;
		data_a[1317]<=8'd220;
		data_a[1318]<=8'd219;
		data_a[1319]<=8'd223;
		data_a[1320]<=8'd221;
		data_a[1321]<=8'd223;
		data_a[1322]<=8'd222;
		data_a[1323]<=8'd222;
		data_a[1324]<=8'd223;
		data_a[1325]<=8'd223;
		data_a[1326]<=8'd221;
		data_a[1327]<=8'd222;
		data_a[1328]<=8'd224;
		data_a[1329]<=8'd229;
		data_a[1330]<=8'd230;
		data_a[1331]<=8'd228;
		data_a[1332]<=8'd231;
		data_a[1333]<=8'd234;
		data_a[1334]<=8'd235;
		data_a[1335]<=8'd240;
		data_a[1336]<=8'd239;
		data_a[1337]<=8'd240;
		data_a[1338]<=8'd243;
		data_a[1339]<=8'd247;
		data_a[1340]<=8'd251;
		data_a[1341]<=8'd253;
		data_a[1342]<=8'd253;
		data_a[1343]<=8'd253;
		data_a[1344]<=8'd255;
		data_a[1345]<=8'd255;
		data_a[1346]<=8'd255;
		data_a[1347]<=8'd255;
		data_a[1348]<=8'd255;
		data_a[1349]<=8'd255;
		data_a[1350]<=8'd255;
		data_a[1351]<=8'd232;
		data_a[1352]<=8'd229;
		data_a[1353]<=8'd231;
		data_a[1354]<=8'd223;
		data_a[1355]<=8'd226;
		data_a[1356]<=8'd223;
		data_a[1357]<=8'd222;
		data_a[1358]<=8'd220;
		data_a[1359]<=8'd220;
		data_a[1360]<=8'd219;
		data_a[1361]<=8'd219;
		data_a[1362]<=8'd219;
		data_a[1363]<=8'd219;
		data_a[1364]<=8'd219;
		data_a[1365]<=8'd219;
		data_a[1366]<=8'd218;
		data_a[1367]<=8'd218;
		data_a[1368]<=8'd217;
		data_a[1369]<=8'd217;
		data_a[1370]<=8'd217;
		data_a[1371]<=8'd217;
		data_a[1372]<=8'd217;
		data_a[1373]<=8'd217;
		data_a[1374]<=8'd218;
		data_a[1375]<=8'd218;
		data_a[1376]<=8'd217;
		data_a[1377]<=8'd215;
		data_a[1378]<=8'd216;
		data_a[1379]<=8'd219;
		data_a[1380]<=8'd219;
		data_a[1381]<=8'd216;
		data_a[1382]<=8'd221;
		data_a[1383]<=8'd216;
		data_a[1384]<=8'd211;
		data_a[1385]<=8'd218;
		data_a[1386]<=8'd218;
		data_a[1387]<=8'd220;
		data_a[1388]<=8'd217;
		data_a[1389]<=8'd220;
		data_a[1390]<=8'd217;
		data_a[1391]<=8'd210;
		data_a[1392]<=8'd210;
		data_a[1393]<=8'd218;
		data_a[1394]<=8'd223;
		data_a[1395]<=8'd222;
		data_a[1396]<=8'd224;
		data_a[1397]<=8'd228;
		data_a[1398]<=8'd227;
		data_a[1399]<=8'd231;
		data_a[1400]<=8'd232;
		data_a[1401]<=8'd238;
		data_a[1402]<=8'd239;
		data_a[1403]<=8'd249;
		data_a[1404]<=8'd253;
		data_a[1405]<=8'd255;
		data_a[1406]<=8'd255;
		data_a[1407]<=8'd255;
		data_a[1408]<=8'd255;
		data_a[1409]<=8'd255;
		data_a[1410]<=8'd254;
		data_a[1411]<=8'd254;
		data_a[1412]<=8'd254;
		data_a[1413]<=8'd253;
		data_a[1414]<=8'd255;
		data_a[1415]<=8'd253;
		data_a[1416]<=8'd249;
		data_a[1417]<=8'd244;
		data_a[1418]<=8'd239;
		data_a[1419]<=8'd236;
		data_a[1420]<=8'd234;
		data_a[1421]<=8'd234;
		data_a[1422]<=8'd227;
		data_a[1423]<=8'd226;
		data_a[1424]<=8'd224;
		data_a[1425]<=8'd222;
		data_a[1426]<=8'd220;
		data_a[1427]<=8'd220;
		data_a[1428]<=8'd220;
		data_a[1429]<=8'd220;
		data_a[1430]<=8'd217;
		data_a[1431]<=8'd220;
		data_a[1432]<=8'd212;
		data_a[1433]<=8'd212;
		data_a[1434]<=8'd218;
		data_a[1435]<=8'd217;
		data_a[1436]<=8'd213;
		data_a[1437]<=8'd215;
		data_a[1438]<=8'd217;
		data_a[1439]<=8'd215;
		data_a[1440]<=8'd214;
		data_a[1441]<=8'd209;
		data_a[1442]<=8'd211;
		data_a[1443]<=8'd217;
		data_a[1444]<=8'd216;
		data_a[1445]<=8'd218;
		data_a[1446]<=8'd215;
		data_a[1447]<=8'd213;
		data_a[1448]<=8'd216;
		data_a[1449]<=8'd218;
		data_a[1450]<=8'd204;
		data_a[1451]<=8'd203;
		data_a[1452]<=8'd209;
		data_a[1453]<=8'd208;
		data_a[1454]<=8'd207;
		data_a[1455]<=8'd191;
		data_a[1456]<=8'd176;
		data_a[1457]<=8'd168;
		data_a[1458]<=8'd167;
		data_a[1459]<=8'd176;
		data_a[1460]<=8'd182;
		data_a[1461]<=8'd145;
		data_a[1462]<=8'd198;
		data_a[1463]<=8'd173;
		data_a[1464]<=8'd208;
		data_a[1465]<=8'd225;
		data_a[1466]<=8'd200;
		data_a[1467]<=8'd221;
		data_a[1468]<=8'd221;
		data_a[1469]<=8'd221;
		data_a[1470]<=8'd218;
		data_a[1471]<=8'd221;
		data_a[1472]<=8'd221;
		data_a[1473]<=8'd221;
		data_a[1474]<=8'd223;
		data_a[1475]<=8'd224;
		data_a[1476]<=8'd223;
		data_a[1477]<=8'd224;
		data_a[1478]<=8'd226;
		data_a[1479]<=8'd229;
		data_a[1480]<=8'd226;
		data_a[1481]<=8'd232;
		data_a[1482]<=8'd238;
		data_a[1483]<=8'd234;
		data_a[1484]<=8'd237;
		data_a[1485]<=8'd239;
		data_a[1486]<=8'd245;
		data_a[1487]<=8'd246;
		data_a[1488]<=8'd249;
		data_a[1489]<=8'd252;
		data_a[1490]<=8'd253;
		data_a[1491]<=8'd254;
		data_a[1492]<=8'd254;
		data_a[1493]<=8'd254;
		data_a[1494]<=8'd255;
		data_a[1495]<=8'd255;
		data_a[1496]<=8'd255;
		data_a[1497]<=8'd255;
		data_a[1498]<=8'd255;
		data_a[1499]<=8'd255;
		data_a[1500]<=8'd253;
		data_a[1501]<=8'd255;
		data_a[1502]<=8'd233;
		data_a[1503]<=8'd230;
		data_a[1504]<=8'd233;
		data_a[1505]<=8'd225;
		data_a[1506]<=8'd222;
		data_a[1507]<=8'd220;
		data_a[1508]<=8'd219;
		data_a[1509]<=8'd219;
		data_a[1510]<=8'd219;
		data_a[1511]<=8'd219;
		data_a[1512]<=8'd219;
		data_a[1513]<=8'd219;
		data_a[1514]<=8'd220;
		data_a[1515]<=8'd220;
		data_a[1516]<=8'd217;
		data_a[1517]<=8'd217;
		data_a[1518]<=8'd217;
		data_a[1519]<=8'd217;
		data_a[1520]<=8'd217;
		data_a[1521]<=8'd216;
		data_a[1522]<=8'd216;
		data_a[1523]<=8'd217;
		data_a[1524]<=8'd214;
		data_a[1525]<=8'd218;
		data_a[1526]<=8'd220;
		data_a[1527]<=8'd217;
		data_a[1528]<=8'd215;
		data_a[1529]<=8'd216;
		data_a[1530]<=8'd218;
		data_a[1531]<=8'd219;
		data_a[1532]<=8'd214;
		data_a[1533]<=8'd217;
		data_a[1534]<=8'd215;
		data_a[1535]<=8'd216;
		data_a[1536]<=8'd212;
		data_a[1537]<=8'd216;
		data_a[1538]<=8'd213;
		data_a[1539]<=8'd212;
		data_a[1540]<=8'd208;
		data_a[1541]<=8'd216;
		data_a[1542]<=8'd222;
		data_a[1543]<=8'd221;
		data_a[1544]<=8'd219;
		data_a[1545]<=8'd221;
		data_a[1546]<=8'd224;
		data_a[1547]<=8'd225;
		data_a[1548]<=8'd227;
		data_a[1549]<=8'd228;
		data_a[1550]<=8'd231;
		data_a[1551]<=8'd238;
		data_a[1552]<=8'd240;
		data_a[1553]<=8'd244;
		data_a[1554]<=8'd248;
		data_a[1555]<=8'd255;
		data_a[1556]<=8'd254;
		data_a[1557]<=8'd254;
		data_a[1558]<=8'd254;
		data_a[1559]<=8'd255;
		data_a[1560]<=8'd255;
		data_a[1561]<=8'd255;
		data_a[1562]<=8'd255;
		data_a[1563]<=8'd255;
		data_a[1564]<=8'd249;
		data_a[1565]<=8'd245;
		data_a[1566]<=8'd240;
		data_a[1567]<=8'd236;
		data_a[1568]<=8'd234;
		data_a[1569]<=8'd233;
		data_a[1570]<=8'd233;
		data_a[1571]<=8'd232;
		data_a[1572]<=8'd227;
		data_a[1573]<=8'd225;
		data_a[1574]<=8'd223;
		data_a[1575]<=8'd222;
		data_a[1576]<=8'd221;
		data_a[1577]<=8'd221;
		data_a[1578]<=8'd220;
		data_a[1579]<=8'd219;
		data_a[1580]<=8'd219;
		data_a[1581]<=8'd219;
		data_a[1582]<=8'd213;
		data_a[1583]<=8'd217;
		data_a[1584]<=8'd218;
		data_a[1585]<=8'd216;
		data_a[1586]<=8'd215;
		data_a[1587]<=8'd215;
		data_a[1588]<=8'd215;
		data_a[1589]<=8'd209;
		data_a[1590]<=8'd214;
		data_a[1591]<=8'd215;
		data_a[1592]<=8'd216;
		data_a[1593]<=8'd207;
		data_a[1594]<=8'd212;
		data_a[1595]<=8'd200;
		data_a[1596]<=8'd188;
		data_a[1597]<=8'd209;
		data_a[1598]<=8'd223;
		data_a[1599]<=8'd218;
		data_a[1600]<=8'd182;
		data_a[1601]<=8'd158;
		data_a[1602]<=8'd159;
		data_a[1603]<=8'd171;
		data_a[1604]<=8'd169;
		data_a[1605]<=8'd167;
		data_a[1606]<=8'd166;
		data_a[1607]<=8'd148;
		data_a[1608]<=8'd138;
		data_a[1609]<=8'd143;
		data_a[1610]<=8'd180;
		data_a[1611]<=8'd167;
		data_a[1612]<=8'd165;
		data_a[1613]<=8'd171;
		data_a[1614]<=8'd199;
		data_a[1615]<=8'd205;
		data_a[1616]<=8'd212;
		data_a[1617]<=8'd218;
		data_a[1618]<=8'd216;
		data_a[1619]<=8'd221;
		data_a[1620]<=8'd218;
		data_a[1621]<=8'd221;
		data_a[1622]<=8'd221;
		data_a[1623]<=8'd220;
		data_a[1624]<=8'd222;
		data_a[1625]<=8'd224;
		data_a[1626]<=8'd223;
		data_a[1627]<=8'd224;
		data_a[1628]<=8'd223;
		data_a[1629]<=8'd228;
		data_a[1630]<=8'd235;
		data_a[1631]<=8'd230;
		data_a[1632]<=8'd233;
		data_a[1633]<=8'd242;
		data_a[1634]<=8'd240;
		data_a[1635]<=8'd246;
		data_a[1636]<=8'd251;
		data_a[1637]<=8'd253;
		data_a[1638]<=8'd254;
		data_a[1639]<=8'd255;
		data_a[1640]<=8'd255;
		data_a[1641]<=8'd255;
		data_a[1642]<=8'd255;
		data_a[1643]<=8'd255;
		data_a[1644]<=8'd254;
		data_a[1645]<=8'd254;
		data_a[1646]<=8'd254;
		data_a[1647]<=8'd254;
		data_a[1648]<=8'd254;
		data_a[1649]<=8'd254;
		data_a[1650]<=8'd255;
		data_a[1651]<=8'd253;
		data_a[1652]<=8'd255;
		data_a[1653]<=8'd244;
		data_a[1654]<=8'd223;
		data_a[1655]<=8'd224;
		data_a[1656]<=8'd217;
		data_a[1657]<=8'd225;
		data_a[1658]<=8'd220;
		data_a[1659]<=8'd220;
		data_a[1660]<=8'd220;
		data_a[1661]<=8'd220;
		data_a[1662]<=8'd219;
		data_a[1663]<=8'd219;
		data_a[1664]<=8'd219;
		data_a[1665]<=8'd219;
		data_a[1666]<=8'd217;
		data_a[1667]<=8'd217;
		data_a[1668]<=8'd218;
		data_a[1669]<=8'd217;
		data_a[1670]<=8'd217;
		data_a[1671]<=8'd216;
		data_a[1672]<=8'd216;
		data_a[1673]<=8'd217;
		data_a[1674]<=8'd220;
		data_a[1675]<=8'd216;
		data_a[1676]<=8'd214;
		data_a[1677]<=8'd216;
		data_a[1678]<=8'd217;
		data_a[1679]<=8'd217;
		data_a[1680]<=8'd218;
		data_a[1681]<=8'd221;
		data_a[1682]<=8'd220;
		data_a[1683]<=8'd214;
		data_a[1684]<=8'd216;
		data_a[1685]<=8'd216;
		data_a[1686]<=8'd217;
		data_a[1687]<=8'd207;
		data_a[1688]<=8'd210;
		data_a[1689]<=8'd216;
		data_a[1690]<=8'd217;
		data_a[1691]<=8'd218;
		data_a[1692]<=8'd220;
		data_a[1693]<=8'd220;
		data_a[1694]<=8'd220;
		data_a[1695]<=8'd221;
		data_a[1696]<=8'd222;
		data_a[1697]<=8'd223;
		data_a[1698]<=8'd228;
		data_a[1699]<=8'd228;
		data_a[1700]<=8'd230;
		data_a[1701]<=8'd235;
		data_a[1702]<=8'd237;
		data_a[1703]<=8'd238;
		data_a[1704]<=8'd241;
		data_a[1705]<=8'd247;
		data_a[1706]<=8'd255;
		data_a[1707]<=8'd255;
		data_a[1708]<=8'd255;
		data_a[1709]<=8'd255;
		data_a[1710]<=8'd252;
		data_a[1711]<=8'd249;
		data_a[1712]<=8'd247;
		data_a[1713]<=8'd246;
		data_a[1714]<=8'd243;
		data_a[1715]<=8'd242;
		data_a[1716]<=8'd240;
		data_a[1717]<=8'd239;
		data_a[1718]<=8'd238;
		data_a[1719]<=8'd236;
		data_a[1720]<=8'd234;
		data_a[1721]<=8'd231;
		data_a[1722]<=8'd227;
		data_a[1723]<=8'd225;
		data_a[1724]<=8'd223;
		data_a[1725]<=8'd222;
		data_a[1726]<=8'd221;
		data_a[1727]<=8'd221;
		data_a[1728]<=8'd219;
		data_a[1729]<=8'd218;
		data_a[1730]<=8'd218;
		data_a[1731]<=8'd219;
		data_a[1732]<=8'd218;
		data_a[1733]<=8'd220;
		data_a[1734]<=8'd213;
		data_a[1735]<=8'd219;
		data_a[1736]<=8'd213;
		data_a[1737]<=8'd212;
		data_a[1738]<=8'd214;
		data_a[1739]<=8'd219;
		data_a[1740]<=8'd218;
		data_a[1741]<=8'd174;
		data_a[1742]<=8'd186;
		data_a[1743]<=8'd149;
		data_a[1744]<=8'd171;
		data_a[1745]<=8'd164;
		data_a[1746]<=8'd119;
		data_a[1747]<=8'd127;
		data_a[1748]<=8'd147;
		data_a[1749]<=8'd175;
		data_a[1750]<=8'd164;
		data_a[1751]<=8'd165;
		data_a[1752]<=8'd169;
		data_a[1753]<=8'd151;
		data_a[1754]<=8'd133;
		data_a[1755]<=8'd160;
		data_a[1756]<=8'd139;
		data_a[1757]<=8'd141;
		data_a[1758]<=8'd153;
		data_a[1759]<=8'd140;
		data_a[1760]<=8'd144;
		data_a[1761]<=8'd162;
		data_a[1762]<=8'd165;
		data_a[1763]<=8'd142;
		data_a[1764]<=8'd172;
		data_a[1765]<=8'd186;
		data_a[1766]<=8'd200;
		data_a[1767]<=8'd202;
		data_a[1768]<=8'd222;
		data_a[1769]<=8'd220;
		data_a[1770]<=8'd219;
		data_a[1771]<=8'd222;
		data_a[1772]<=8'd221;
		data_a[1773]<=8'd219;
		data_a[1774]<=8'd222;
		data_a[1775]<=8'd223;
		data_a[1776]<=8'd222;
		data_a[1777]<=8'd223;
		data_a[1778]<=8'd225;
		data_a[1779]<=8'd226;
		data_a[1780]<=8'd224;
		data_a[1781]<=8'd236;
		data_a[1782]<=8'd240;
		data_a[1783]<=8'd236;
		data_a[1784]<=8'd249;
		data_a[1785]<=8'd255;
		data_a[1786]<=8'd255;
		data_a[1787]<=8'd255;
		data_a[1788]<=8'd255;
		data_a[1789]<=8'd255;
		data_a[1790]<=8'd255;
		data_a[1791]<=8'd255;
		data_a[1792]<=8'd255;
		data_a[1793]<=8'd255;
		data_a[1794]<=8'd254;
		data_a[1795]<=8'd254;
		data_a[1796]<=8'd254;
		data_a[1797]<=8'd254;
		data_a[1798]<=8'd254;
		data_a[1799]<=8'd254;
		data_a[1800]<=8'd254;
		data_a[1801]<=8'd255;
		data_a[1802]<=8'd253;
		data_a[1803]<=8'd254;
		data_a[1804]<=8'd223;
		data_a[1805]<=8'd228;
		data_a[1806]<=8'd220;
		data_a[1807]<=8'd226;
		data_a[1808]<=8'd219;
		data_a[1809]<=8'd219;
		data_a[1810]<=8'd219;
		data_a[1811]<=8'd219;
		data_a[1812]<=8'd219;
		data_a[1813]<=8'd218;
		data_a[1814]<=8'd218;
		data_a[1815]<=8'd218;
		data_a[1816]<=8'd217;
		data_a[1817]<=8'd217;
		data_a[1818]<=8'd217;
		data_a[1819]<=8'd217;
		data_a[1820]<=8'd217;
		data_a[1821]<=8'd216;
		data_a[1822]<=8'd216;
		data_a[1823]<=8'd216;
		data_a[1824]<=8'd221;
		data_a[1825]<=8'd217;
		data_a[1826]<=8'd215;
		data_a[1827]<=8'd216;
		data_a[1828]<=8'd215;
		data_a[1829]<=8'd214;
		data_a[1830]<=8'd218;
		data_a[1831]<=8'd225;
		data_a[1832]<=8'd216;
		data_a[1833]<=8'd216;
		data_a[1834]<=8'd214;
		data_a[1835]<=8'd205;
		data_a[1836]<=8'd210;
		data_a[1837]<=8'd216;
		data_a[1838]<=8'd221;
		data_a[1839]<=8'd215;
		data_a[1840]<=8'd217;
		data_a[1841]<=8'd217;
		data_a[1842]<=8'd217;
		data_a[1843]<=8'd217;
		data_a[1844]<=8'd218;
		data_a[1845]<=8'd221;
		data_a[1846]<=8'd224;
		data_a[1847]<=8'd226;
		data_a[1848]<=8'd228;
		data_a[1849]<=8'd227;
		data_a[1850]<=8'd229;
		data_a[1851]<=8'd231;
		data_a[1852]<=8'd234;
		data_a[1853]<=8'd234;
		data_a[1854]<=8'd237;
		data_a[1855]<=8'd239;
		data_a[1856]<=8'd249;
		data_a[1857]<=8'd252;
		data_a[1858]<=8'd254;
		data_a[1859]<=8'd253;
		data_a[1860]<=8'd248;
		data_a[1861]<=8'd243;
		data_a[1862]<=8'd242;
		data_a[1863]<=8'd242;
		data_a[1864]<=8'd239;
		data_a[1865]<=8'd240;
		data_a[1866]<=8'd240;
		data_a[1867]<=8'd240;
		data_a[1868]<=8'd238;
		data_a[1869]<=8'd234;
		data_a[1870]<=8'd230;
		data_a[1871]<=8'd227;
		data_a[1872]<=8'd226;
		data_a[1873]<=8'd225;
		data_a[1874]<=8'd223;
		data_a[1875]<=8'd221;
		data_a[1876]<=8'd220;
		data_a[1877]<=8'd220;
		data_a[1878]<=8'd219;
		data_a[1879]<=8'd219;
		data_a[1880]<=8'd216;
		data_a[1881]<=8'd219;
		data_a[1882]<=8'd217;
		data_a[1883]<=8'd214;
		data_a[1884]<=8'd211;
		data_a[1885]<=8'd214;
		data_a[1886]<=8'd216;
		data_a[1887]<=8'd210;
		data_a[1888]<=8'd203;
		data_a[1889]<=8'd206;
		data_a[1890]<=8'd178;
		data_a[1891]<=8'd158;
		data_a[1892]<=8'd150;
		data_a[1893]<=8'd165;
		data_a[1894]<=8'd175;
		data_a[1895]<=8'd158;
		data_a[1896]<=8'd144;
		data_a[1897]<=8'd116;
		data_a[1898]<=8'd94;
		data_a[1899]<=8'd129;
		data_a[1900]<=8'd155;
		data_a[1901]<=8'd159;
		data_a[1902]<=8'd163;
		data_a[1903]<=8'd157;
		data_a[1904]<=8'd153;
		data_a[1905]<=8'd134;
		data_a[1906]<=8'd140;
		data_a[1907]<=8'd144;
		data_a[1908]<=8'd141;
		data_a[1909]<=8'd124;
		data_a[1910]<=8'd115;
		data_a[1911]<=8'd133;
		data_a[1912]<=8'd154;
		data_a[1913]<=8'd166;
		data_a[1914]<=8'd146;
		data_a[1915]<=8'd177;
		data_a[1916]<=8'd178;
		data_a[1917]<=8'd194;
		data_a[1918]<=8'd217;
		data_a[1919]<=8'd216;
		data_a[1920]<=8'd218;
		data_a[1921]<=8'd221;
		data_a[1922]<=8'd220;
		data_a[1923]<=8'd218;
		data_a[1924]<=8'd221;
		data_a[1925]<=8'd223;
		data_a[1926]<=8'd223;
		data_a[1927]<=8'd223;
		data_a[1928]<=8'd225;
		data_a[1929]<=8'd222;
		data_a[1930]<=8'd231;
		data_a[1931]<=8'd232;
		data_a[1932]<=8'd243;
		data_a[1933]<=8'd255;
		data_a[1934]<=8'd254;
		data_a[1935]<=8'd254;
		data_a[1936]<=8'd255;
		data_a[1937]<=8'd255;
		data_a[1938]<=8'd254;
		data_a[1939]<=8'd254;
		data_a[1940]<=8'd255;
		data_a[1941]<=8'd255;
		data_a[1942]<=8'd254;
		data_a[1943]<=8'd254;
		data_a[1944]<=8'd254;
		data_a[1945]<=8'd254;
		data_a[1946]<=8'd254;
		data_a[1947]<=8'd254;
		data_a[1948]<=8'd254;
		data_a[1949]<=8'd254;
		data_a[1950]<=8'd254;
		data_a[1951]<=8'd255;
		data_a[1952]<=8'd255;
		data_a[1953]<=8'd254;
		data_a[1954]<=8'd252;
		data_a[1955]<=8'd198;
		data_a[1956]<=8'd214;
		data_a[1957]<=8'd223;
		data_a[1958]<=8'd219;
		data_a[1959]<=8'd219;
		data_a[1960]<=8'd219;
		data_a[1961]<=8'd219;
		data_a[1962]<=8'd218;
		data_a[1963]<=8'd219;
		data_a[1964]<=8'd219;
		data_a[1965]<=8'd219;
		data_a[1966]<=8'd217;
		data_a[1967]<=8'd217;
		data_a[1968]<=8'd216;
		data_a[1969]<=8'd216;
		data_a[1970]<=8'd216;
		data_a[1971]<=8'd216;
		data_a[1972]<=8'd216;
		data_a[1973]<=8'd215;
		data_a[1974]<=8'd215;
		data_a[1975]<=8'd217;
		data_a[1976]<=8'd218;
		data_a[1977]<=8'd217;
		data_a[1978]<=8'd216;
		data_a[1979]<=8'd216;
		data_a[1980]<=8'd216;
		data_a[1981]<=8'd216;
		data_a[1982]<=8'd210;
		data_a[1983]<=8'd210;
		data_a[1984]<=8'd207;
		data_a[1985]<=8'd212;
		data_a[1986]<=8'd211;
		data_a[1987]<=8'd215;
		data_a[1988]<=8'd215;
		data_a[1989]<=8'd219;
		data_a[1990]<=8'd214;
		data_a[1991]<=8'd218;
		data_a[1992]<=8'd220;
		data_a[1993]<=8'd217;
		data_a[1994]<=8'd215;
		data_a[1995]<=8'd218;
		data_a[1996]<=8'd222;
		data_a[1997]<=8'd225;
		data_a[1998]<=8'd226;
		data_a[1999]<=8'd227;
		data_a[2000]<=8'd230;
		data_a[2001]<=8'd230;
		data_a[2002]<=8'd234;
		data_a[2003]<=8'd235;
		data_a[2004]<=8'd239;
		data_a[2005]<=8'd238;
		data_a[2006]<=8'd229;
		data_a[2007]<=8'd234;
		data_a[2008]<=8'd239;
		data_a[2009]<=8'd241;
		data_a[2010]<=8'd239;
		data_a[2011]<=8'd237;
		data_a[2012]<=8'd238;
		data_a[2013]<=8'd240;
		data_a[2014]<=8'd236;
		data_a[2015]<=8'd237;
		data_a[2016]<=8'd236;
		data_a[2017]<=8'd235;
		data_a[2018]<=8'd233;
		data_a[2019]<=8'd230;
		data_a[2020]<=8'd228;
		data_a[2021]<=8'd227;
		data_a[2022]<=8'd225;
		data_a[2023]<=8'd224;
		data_a[2024]<=8'd223;
		data_a[2025]<=8'd221;
		data_a[2026]<=8'd220;
		data_a[2027]<=8'd219;
		data_a[2028]<=8'd218;
		data_a[2029]<=8'd218;
		data_a[2030]<=8'd219;
		data_a[2031]<=8'd212;
		data_a[2032]<=8'd220;
		data_a[2033]<=8'd210;
		data_a[2034]<=8'd218;
		data_a[2035]<=8'd215;
		data_a[2036]<=8'd214;
		data_a[2037]<=8'd228;
		data_a[2038]<=8'd143;
		data_a[2039]<=8'd144;
		data_a[2040]<=8'd144;
		data_a[2041]<=8'd143;
		data_a[2042]<=8'd140;
		data_a[2043]<=8'd152;
		data_a[2044]<=8'd163;
		data_a[2045]<=8'd149;
		data_a[2046]<=8'd148;
		data_a[2047]<=8'd125;
		data_a[2048]<=8'd116;
		data_a[2049]<=8'd122;
		data_a[2050]<=8'd121;
		data_a[2051]<=8'd131;
		data_a[2052]<=8'd154;
		data_a[2053]<=8'd153;
		data_a[2054]<=8'd145;
		data_a[2055]<=8'd151;
		data_a[2056]<=8'd150;
		data_a[2057]<=8'd152;
		data_a[2058]<=8'd132;
		data_a[2059]<=8'd152;
		data_a[2060]<=8'd128;
		data_a[2061]<=8'd127;
		data_a[2062]<=8'd124;
		data_a[2063]<=8'd167;
		data_a[2064]<=8'd141;
		data_a[2065]<=8'd160;
		data_a[2066]<=8'd171;
		data_a[2067]<=8'd202;
		data_a[2068]<=8'd190;
		data_a[2069]<=8'd219;
		data_a[2070]<=8'd218;
		data_a[2071]<=8'd221;
		data_a[2072]<=8'd220;
		data_a[2073]<=8'd217;
		data_a[2074]<=8'd219;
		data_a[2075]<=8'd222;
		data_a[2076]<=8'd222;
		data_a[2077]<=8'd222;
		data_a[2078]<=8'd225;
		data_a[2079]<=8'd223;
		data_a[2080]<=8'd228;
		data_a[2081]<=8'd249;
		data_a[2082]<=8'd255;
		data_a[2083]<=8'd253;
		data_a[2084]<=8'd255;
		data_a[2085]<=8'd254;
		data_a[2086]<=8'd255;
		data_a[2087]<=8'd255;
		data_a[2088]<=8'd254;
		data_a[2089]<=8'd254;
		data_a[2090]<=8'd254;
		data_a[2091]<=8'd254;
		data_a[2092]<=8'd254;
		data_a[2093]<=8'd254;
		data_a[2094]<=8'd255;
		data_a[2095]<=8'd255;
		data_a[2096]<=8'd255;
		data_a[2097]<=8'd255;
		data_a[2098]<=8'd255;
		data_a[2099]<=8'd255;
		data_a[2100]<=8'd254;
		data_a[2101]<=8'd254;
		data_a[2102]<=8'd255;
		data_a[2103]<=8'd255;
		data_a[2104]<=8'd253;
		data_a[2105]<=8'd255;
		data_a[2106]<=8'd228;
		data_a[2107]<=8'd217;
		data_a[2108]<=8'd220;
		data_a[2109]<=8'd220;
		data_a[2110]<=8'd219;
		data_a[2111]<=8'd218;
		data_a[2112]<=8'd218;
		data_a[2113]<=8'd218;
		data_a[2114]<=8'd218;
		data_a[2115]<=8'd218;
		data_a[2116]<=8'd217;
		data_a[2117]<=8'd216;
		data_a[2118]<=8'd215;
		data_a[2119]<=8'd215;
		data_a[2120]<=8'd216;
		data_a[2121]<=8'd216;
		data_a[2122]<=8'd215;
		data_a[2123]<=8'd214;
		data_a[2124]<=8'd217;
		data_a[2125]<=8'd214;
		data_a[2126]<=8'd213;
		data_a[2127]<=8'd215;
		data_a[2128]<=8'd218;
		data_a[2129]<=8'd218;
		data_a[2130]<=8'd213;
		data_a[2131]<=8'd206;
		data_a[2132]<=8'd208;
		data_a[2133]<=8'd216;
		data_a[2134]<=8'd217;
		data_a[2135]<=8'd218;
		data_a[2136]<=8'd213;
		data_a[2137]<=8'd217;
		data_a[2138]<=8'd216;
		data_a[2139]<=8'd216;
		data_a[2140]<=8'd222;
		data_a[2141]<=8'd213;
		data_a[2142]<=8'd212;
		data_a[2143]<=8'd220;
		data_a[2144]<=8'd222;
		data_a[2145]<=8'd217;
		data_a[2146]<=8'd216;
		data_a[2147]<=8'd222;
		data_a[2148]<=8'd225;
		data_a[2149]<=8'd226;
		data_a[2150]<=8'd230;
		data_a[2151]<=8'd230;
		data_a[2152]<=8'd235;
		data_a[2153]<=8'd234;
		data_a[2154]<=8'd239;
		data_a[2155]<=8'd239;
		data_a[2156]<=8'd235;
		data_a[2157]<=8'd238;
		data_a[2158]<=8'd240;
		data_a[2159]<=8'd241;
		data_a[2160]<=8'd241;
		data_a[2161]<=8'd240;
		data_a[2162]<=8'd240;
		data_a[2163]<=8'd241;
		data_a[2164]<=8'd237;
		data_a[2165]<=8'd237;
		data_a[2166]<=8'd236;
		data_a[2167]<=8'd234;
		data_a[2168]<=8'd232;
		data_a[2169]<=8'd231;
		data_a[2170]<=8'd231;
		data_a[2171]<=8'd231;
		data_a[2172]<=8'd223;
		data_a[2173]<=8'd224;
		data_a[2174]<=8'd223;
		data_a[2175]<=8'd222;
		data_a[2176]<=8'd219;
		data_a[2177]<=8'd218;
		data_a[2178]<=8'd217;
		data_a[2179]<=8'd218;
		data_a[2180]<=8'd214;
		data_a[2181]<=8'd219;
		data_a[2182]<=8'd213;
		data_a[2183]<=8'd217;
		data_a[2184]<=8'd214;
		data_a[2185]<=8'd216;
		data_a[2186]<=8'd196;
		data_a[2187]<=8'd117;
		data_a[2188]<=8'd145;
		data_a[2189]<=8'd151;
		data_a[2190]<=8'd148;
		data_a[2191]<=8'd146;
		data_a[2192]<=8'd160;
		data_a[2193]<=8'd153;
		data_a[2194]<=8'd134;
		data_a[2195]<=8'd138;
		data_a[2196]<=8'd133;
		data_a[2197]<=8'd115;
		data_a[2198]<=8'd129;
		data_a[2199]<=8'd134;
		data_a[2200]<=8'd132;
		data_a[2201]<=8'd116;
		data_a[2202]<=8'd116;
		data_a[2203]<=8'd140;
		data_a[2204]<=8'd155;
		data_a[2205]<=8'd158;
		data_a[2206]<=8'd154;
		data_a[2207]<=8'd156;
		data_a[2208]<=8'd149;
		data_a[2209]<=8'd120;
		data_a[2210]<=8'd133;
		data_a[2211]<=8'd126;
		data_a[2212]<=8'd128;
		data_a[2213]<=8'd133;
		data_a[2214]<=8'd144;
		data_a[2215]<=8'd120;
		data_a[2216]<=8'd209;
		data_a[2217]<=8'd166;
		data_a[2218]<=8'd206;
		data_a[2219]<=8'd214;
		data_a[2220]<=8'd217;
		data_a[2221]<=8'd220;
		data_a[2222]<=8'd218;
		data_a[2223]<=8'd215;
		data_a[2224]<=8'd217;
		data_a[2225]<=8'd220;
		data_a[2226]<=8'd221;
		data_a[2227]<=8'd220;
		data_a[2228]<=8'd221;
		data_a[2229]<=8'd224;
		data_a[2230]<=8'd242;
		data_a[2231]<=8'd252;
		data_a[2232]<=8'd254;
		data_a[2233]<=8'd255;
		data_a[2234]<=8'd254;
		data_a[2235]<=8'd254;
		data_a[2236]<=8'd255;
		data_a[2237]<=8'd254;
		data_a[2238]<=8'd254;
		data_a[2239]<=8'd254;
		data_a[2240]<=8'd254;
		data_a[2241]<=8'd254;
		data_a[2242]<=8'd254;
		data_a[2243]<=8'd254;
		data_a[2244]<=8'd255;
		data_a[2245]<=8'd255;
		data_a[2246]<=8'd255;
		data_a[2247]<=8'd255;
		data_a[2248]<=8'd255;
		data_a[2249]<=8'd255;
		data_a[2250]<=8'd254;
		data_a[2251]<=8'd254;
		data_a[2252]<=8'd255;
		data_a[2253]<=8'd254;
		data_a[2254]<=8'd255;
		data_a[2255]<=8'd234;
		data_a[2256]<=8'd182;
		data_a[2257]<=8'd201;
		data_a[2258]<=8'd221;
		data_a[2259]<=8'd220;
		data_a[2260]<=8'd218;
		data_a[2261]<=8'd217;
		data_a[2262]<=8'd216;
		data_a[2263]<=8'd216;
		data_a[2264]<=8'd216;
		data_a[2265]<=8'd216;
		data_a[2266]<=8'd216;
		data_a[2267]<=8'd215;
		data_a[2268]<=8'd213;
		data_a[2269]<=8'd214;
		data_a[2270]<=8'd215;
		data_a[2271]<=8'd216;
		data_a[2272]<=8'd215;
		data_a[2273]<=8'd213;
		data_a[2274]<=8'd214;
		data_a[2275]<=8'd215;
		data_a[2276]<=8'd218;
		data_a[2277]<=8'd216;
		data_a[2278]<=8'd207;
		data_a[2279]<=8'd201;
		data_a[2280]<=8'd208;
		data_a[2281]<=8'd220;
		data_a[2282]<=8'd220;
		data_a[2283]<=8'd215;
		data_a[2284]<=8'd216;
		data_a[2285]<=8'd215;
		data_a[2286]<=8'd219;
		data_a[2287]<=8'd214;
		data_a[2288]<=8'd216;
		data_a[2289]<=8'd217;
		data_a[2290]<=8'd211;
		data_a[2291]<=8'd216;
		data_a[2292]<=8'd219;
		data_a[2293]<=8'd217;
		data_a[2294]<=8'd216;
		data_a[2295]<=8'd220;
		data_a[2296]<=8'd222;
		data_a[2297]<=8'd223;
		data_a[2298]<=8'd224;
		data_a[2299]<=8'd224;
		data_a[2300]<=8'd229;
		data_a[2301]<=8'd229;
		data_a[2302]<=8'd233;
		data_a[2303]<=8'd230;
		data_a[2304]<=8'd235;
		data_a[2305]<=8'd237;
		data_a[2306]<=8'd238;
		data_a[2307]<=8'd238;
		data_a[2308]<=8'd237;
		data_a[2309]<=8'd238;
		data_a[2310]<=8'd238;
		data_a[2311]<=8'd238;
		data_a[2312]<=8'd237;
		data_a[2313]<=8'd236;
		data_a[2314]<=8'd236;
		data_a[2315]<=8'd235;
		data_a[2316]<=8'd233;
		data_a[2317]<=8'd232;
		data_a[2318]<=8'd229;
		data_a[2319]<=8'd228;
		data_a[2320]<=8'd226;
		data_a[2321]<=8'd226;
		data_a[2322]<=8'd222;
		data_a[2323]<=8'd223;
		data_a[2324]<=8'd224;
		data_a[2325]<=8'd222;
		data_a[2326]<=8'd220;
		data_a[2327]<=8'd217;
		data_a[2328]<=8'd217;
		data_a[2329]<=8'd217;
		data_a[2330]<=8'd214;
		data_a[2331]<=8'd216;
		data_a[2332]<=8'd215;
		data_a[2333]<=8'd212;
		data_a[2334]<=8'd222;
		data_a[2335]<=8'd197;
		data_a[2336]<=8'd111;
		data_a[2337]<=8'd165;
		data_a[2338]<=8'd128;
		data_a[2339]<=8'd122;
		data_a[2340]<=8'd144;
		data_a[2341]<=8'd134;
		data_a[2342]<=8'd140;
		data_a[2343]<=8'd140;
		data_a[2344]<=8'd133;
		data_a[2345]<=8'd117;
		data_a[2346]<=8'd119;
		data_a[2347]<=8'd97;
		data_a[2348]<=8'd116;
		data_a[2349]<=8'd101;
		data_a[2350]<=8'd112;
		data_a[2351]<=8'd125;
		data_a[2352]<=8'd114;
		data_a[2353]<=8'd117;
		data_a[2354]<=8'd117;
		data_a[2355]<=8'd120;
		data_a[2356]<=8'd126;
		data_a[2357]<=8'd126;
		data_a[2358]<=8'd134;
		data_a[2359]<=8'd144;
		data_a[2360]<=8'd114;
		data_a[2361]<=8'd131;
		data_a[2362]<=8'd113;
		data_a[2363]<=8'd132;
		data_a[2364]<=8'd141;
		data_a[2365]<=8'd116;
		data_a[2366]<=8'd141;
		data_a[2367]<=8'd158;
		data_a[2368]<=8'd198;
		data_a[2369]<=8'd161;
		data_a[2370]<=8'd213;
		data_a[2371]<=8'd217;
		data_a[2372]<=8'd216;
		data_a[2373]<=8'd214;
		data_a[2374]<=8'd217;
		data_a[2375]<=8'd221;
		data_a[2376]<=8'd222;
		data_a[2377]<=8'd222;
		data_a[2378]<=8'd225;
		data_a[2379]<=8'd225;
		data_a[2380]<=8'd237;
		data_a[2381]<=8'd253;
		data_a[2382]<=8'd255;
		data_a[2383]<=8'd254;
		data_a[2384]<=8'd255;
		data_a[2385]<=8'd255;
		data_a[2386]<=8'd254;
		data_a[2387]<=8'd254;
		data_a[2388]<=8'd254;
		data_a[2389]<=8'd254;
		data_a[2390]<=8'd254;
		data_a[2391]<=8'd254;
		data_a[2392]<=8'd254;
		data_a[2393]<=8'd254;
		data_a[2394]<=8'd255;
		data_a[2395]<=8'd255;
		data_a[2396]<=8'd255;
		data_a[2397]<=8'd255;
		data_a[2398]<=8'd255;
		data_a[2399]<=8'd255;
		data_a[2400]<=8'd254;
		data_a[2401]<=8'd253;
		data_a[2402]<=8'd254;
		data_a[2403]<=8'd254;
		data_a[2404]<=8'd203;
		data_a[2405]<=8'd224;
		data_a[2406]<=8'd223;
		data_a[2407]<=8'd221;
		data_a[2408]<=8'd214;
		data_a[2409]<=8'd210;
		data_a[2410]<=8'd215;
		data_a[2411]<=8'd213;
		data_a[2412]<=8'd219;
		data_a[2413]<=8'd215;
		data_a[2414]<=8'd216;
		data_a[2415]<=8'd216;
		data_a[2416]<=8'd217;
		data_a[2417]<=8'd216;
		data_a[2418]<=8'd214;
		data_a[2419]<=8'd213;
		data_a[2420]<=8'd219;
		data_a[2421]<=8'd211;
		data_a[2422]<=8'd210;
		data_a[2423]<=8'd218;
		data_a[2424]<=8'd219;
		data_a[2425]<=8'd216;
		data_a[2426]<=8'd212;
		data_a[2427]<=8'd198;
		data_a[2428]<=8'd206;
		data_a[2429]<=8'd220;
		data_a[2430]<=8'd214;
		data_a[2431]<=8'd220;
		data_a[2432]<=8'd216;
		data_a[2433]<=8'd215;
		data_a[2434]<=8'd215;
		data_a[2435]<=8'd215;
		data_a[2436]<=8'd215;
		data_a[2437]<=8'd214;
		data_a[2438]<=8'd214;
		data_a[2439]<=8'd215;
		data_a[2440]<=8'd217;
		data_a[2441]<=8'd222;
		data_a[2442]<=8'd216;
		data_a[2443]<=8'd219;
		data_a[2444]<=8'd217;
		data_a[2445]<=8'd216;
		data_a[2446]<=8'd221;
		data_a[2447]<=8'd224;
		data_a[2448]<=8'd224;
		data_a[2449]<=8'd222;
		data_a[2450]<=8'd227;
		data_a[2451]<=8'd227;
		data_a[2452]<=8'd228;
		data_a[2453]<=8'd232;
		data_a[2454]<=8'd231;
		data_a[2455]<=8'd234;
		data_a[2456]<=8'd235;
		data_a[2457]<=8'd239;
		data_a[2458]<=8'd231;
		data_a[2459]<=8'd234;
		data_a[2460]<=8'd239;
		data_a[2461]<=8'd237;
		data_a[2462]<=8'd237;
		data_a[2463]<=8'd233;
		data_a[2464]<=8'd233;
		data_a[2465]<=8'd234;
		data_a[2466]<=8'd234;
		data_a[2467]<=8'd232;
		data_a[2468]<=8'd229;
		data_a[2469]<=8'd228;
		data_a[2470]<=8'd226;
		data_a[2471]<=8'd225;
		data_a[2472]<=8'd222;
		data_a[2473]<=8'd223;
		data_a[2474]<=8'd223;
		data_a[2475]<=8'd221;
		data_a[2476]<=8'd219;
		data_a[2477]<=8'd217;
		data_a[2478]<=8'd217;
		data_a[2479]<=8'd218;
		data_a[2480]<=8'd214;
		data_a[2481]<=8'd216;
		data_a[2482]<=8'd218;
		data_a[2483]<=8'd215;
		data_a[2484]<=8'd224;
		data_a[2485]<=8'd106;
		data_a[2486]<=8'd131;
		data_a[2487]<=8'd149;
		data_a[2488]<=8'd99;
		data_a[2489]<=8'd99;
		data_a[2490]<=8'd112;
		data_a[2491]<=8'd121;
		data_a[2492]<=8'd135;
		data_a[2493]<=8'd132;
		data_a[2494]<=8'd119;
		data_a[2495]<=8'd113;
		data_a[2496]<=8'd106;
		data_a[2497]<=8'd110;
		data_a[2498]<=8'd87;
		data_a[2499]<=8'd108;
		data_a[2500]<=8'd104;
		data_a[2501]<=8'd110;
		data_a[2502]<=8'd133;
		data_a[2503]<=8'd120;
		data_a[2504]<=8'd120;
		data_a[2505]<=8'd121;
		data_a[2506]<=8'd119;
		data_a[2507]<=8'd130;
		data_a[2508]<=8'd130;
		data_a[2509]<=8'd129;
		data_a[2510]<=8'd148;
		data_a[2511]<=8'd151;
		data_a[2512]<=8'd113;
		data_a[2513]<=8'd116;
		data_a[2514]<=8'd133;
		data_a[2515]<=8'd121;
		data_a[2516]<=8'd132;
		data_a[2517]<=8'd169;
		data_a[2518]<=8'd165;
		data_a[2519]<=8'd171;
		data_a[2520]<=8'd197;
		data_a[2521]<=8'd195;
		data_a[2522]<=8'd216;
		data_a[2523]<=8'd224;
		data_a[2524]<=8'd218;
		data_a[2525]<=8'd223;
		data_a[2526]<=8'd226;
		data_a[2527]<=8'd221;
		data_a[2528]<=8'd226;
		data_a[2529]<=8'd223;
		data_a[2530]<=8'd226;
		data_a[2531]<=8'd255;
		data_a[2532]<=8'd253;
		data_a[2533]<=8'd253;
		data_a[2534]<=8'd255;
		data_a[2535]<=8'd254;
		data_a[2536]<=8'd254;
		data_a[2537]<=8'd254;
		data_a[2538]<=8'd254;
		data_a[2539]<=8'd254;
		data_a[2540]<=8'd255;
		data_a[2541]<=8'd255;
		data_a[2542]<=8'd255;
		data_a[2543]<=8'd255;
		data_a[2544]<=8'd255;
		data_a[2545]<=8'd254;
		data_a[2546]<=8'd254;
		data_a[2547]<=8'd254;
		data_a[2548]<=8'd254;
		data_a[2549]<=8'd255;
		data_a[2550]<=8'd254;
		data_a[2551]<=8'd254;
		data_a[2552]<=8'd204;
		data_a[2553]<=8'd222;
		data_a[2554]<=8'd228;
		data_a[2555]<=8'd218;
		data_a[2556]<=8'd219;
		data_a[2557]<=8'd218;
		data_a[2558]<=8'd220;
		data_a[2559]<=8'd209;
		data_a[2560]<=8'd207;
		data_a[2561]<=8'd221;
		data_a[2562]<=8'd218;
		data_a[2563]<=8'd214;
		data_a[2564]<=8'd217;
		data_a[2565]<=8'd216;
		data_a[2566]<=8'd216;
		data_a[2567]<=8'd214;
		data_a[2568]<=8'd217;
		data_a[2569]<=8'd216;
		data_a[2570]<=8'd215;
		data_a[2571]<=8'd214;
		data_a[2572]<=8'd219;
		data_a[2573]<=8'd212;
		data_a[2574]<=8'd210;
		data_a[2575]<=8'd191;
		data_a[2576]<=8'd205;
		data_a[2577]<=8'd222;
		data_a[2578]<=8'd211;
		data_a[2579]<=8'd213;
		data_a[2580]<=8'd221;
		data_a[2581]<=8'd212;
		data_a[2582]<=8'd215;
		data_a[2583]<=8'd215;
		data_a[2584]<=8'd215;
		data_a[2585]<=8'd216;
		data_a[2586]<=8'd215;
		data_a[2587]<=8'd214;
		data_a[2588]<=8'd214;
		data_a[2589]<=8'd214;
		data_a[2590]<=8'd214;
		data_a[2591]<=8'd214;
		data_a[2592]<=8'd217;
		data_a[2593]<=8'd213;
		data_a[2594]<=8'd219;
		data_a[2595]<=8'd217;
		data_a[2596]<=8'd219;
		data_a[2597]<=8'd219;
		data_a[2598]<=8'd222;
		data_a[2599]<=8'd221;
		data_a[2600]<=8'd227;
		data_a[2601]<=8'd227;
		data_a[2602]<=8'd229;
		data_a[2603]<=8'd232;
		data_a[2604]<=8'd231;
		data_a[2605]<=8'd235;
		data_a[2606]<=8'd236;
		data_a[2607]<=8'd236;
		data_a[2608]<=8'd233;
		data_a[2609]<=8'd230;
		data_a[2610]<=8'd232;
		data_a[2611]<=8'd236;
		data_a[2612]<=8'd235;
		data_a[2613]<=8'd234;
		data_a[2614]<=8'd234;
		data_a[2615]<=8'd234;
		data_a[2616]<=8'd233;
		data_a[2617]<=8'd231;
		data_a[2618]<=8'd228;
		data_a[2619]<=8'd227;
		data_a[2620]<=8'd225;
		data_a[2621]<=8'd223;
		data_a[2622]<=8'd222;
		data_a[2623]<=8'd222;
		data_a[2624]<=8'd220;
		data_a[2625]<=8'd219;
		data_a[2626]<=8'd217;
		data_a[2627]<=8'd217;
		data_a[2628]<=8'd217;
		data_a[2629]<=8'd217;
		data_a[2630]<=8'd215;
		data_a[2631]<=8'd213;
		data_a[2632]<=8'd213;
		data_a[2633]<=8'd215;
		data_a[2634]<=8'd151;
		data_a[2635]<=8'd149;
		data_a[2636]<=8'd144;
		data_a[2637]<=8'd132;
		data_a[2638]<=8'd107;
		data_a[2639]<=8'd95;
		data_a[2640]<=8'd93;
		data_a[2641]<=8'd100;
		data_a[2642]<=8'd102;
		data_a[2643]<=8'd113;
		data_a[2644]<=8'd114;
		data_a[2645]<=8'd116;
		data_a[2646]<=8'd110;
		data_a[2647]<=8'd100;
		data_a[2648]<=8'd116;
		data_a[2649]<=8'd143;
		data_a[2650]<=8'd127;
		data_a[2651]<=8'd118;
		data_a[2652]<=8'd118;
		data_a[2653]<=8'd115;
		data_a[2654]<=8'd115;
		data_a[2655]<=8'd125;
		data_a[2656]<=8'd136;
		data_a[2657]<=8'd136;
		data_a[2658]<=8'd129;
		data_a[2659]<=8'd127;
		data_a[2660]<=8'd129;
		data_a[2661]<=8'd126;
		data_a[2662]<=8'd124;
		data_a[2663]<=8'd113;
		data_a[2664]<=8'd116;
		data_a[2665]<=8'd122;
		data_a[2666]<=8'd140;
		data_a[2667]<=8'd141;
		data_a[2668]<=8'd155;
		data_a[2669]<=8'd158;
		data_a[2670]<=8'd166;
		data_a[2671]<=8'd196;
		data_a[2672]<=8'd219;
		data_a[2673]<=8'd221;
		data_a[2674]<=8'd219;
		data_a[2675]<=8'd225;
		data_a[2676]<=8'd221;
		data_a[2677]<=8'd225;
		data_a[2678]<=8'd223;
		data_a[2679]<=8'd226;
		data_a[2680]<=8'd229;
		data_a[2681]<=8'd255;
		data_a[2682]<=8'd253;
		data_a[2683]<=8'd255;
		data_a[2684]<=8'd255;
		data_a[2685]<=8'd255;
		data_a[2686]<=8'd254;
		data_a[2687]<=8'd254;
		data_a[2688]<=8'd254;
		data_a[2689]<=8'd255;
		data_a[2690]<=8'd255;
		data_a[2691]<=8'd255;
		data_a[2692]<=8'd255;
		data_a[2693]<=8'd255;
		data_a[2694]<=8'd255;
		data_a[2695]<=8'd255;
		data_a[2696]<=8'd255;
		data_a[2697]<=8'd255;
		data_a[2698]<=8'd255;
		data_a[2699]<=8'd255;
		data_a[2700]<=8'd250;
		data_a[2701]<=8'd228;
		data_a[2702]<=8'd225;
		data_a[2703]<=8'd235;
		data_a[2704]<=8'd219;
		data_a[2705]<=8'd221;
		data_a[2706]<=8'd213;
		data_a[2707]<=8'd222;
		data_a[2708]<=8'd220;
		data_a[2709]<=8'd211;
		data_a[2710]<=8'd210;
		data_a[2711]<=8'd208;
		data_a[2712]<=8'd217;
		data_a[2713]<=8'd217;
		data_a[2714]<=8'd218;
		data_a[2715]<=8'd217;
		data_a[2716]<=8'd215;
		data_a[2717]<=8'd218;
		data_a[2718]<=8'd216;
		data_a[2719]<=8'd214;
		data_a[2720]<=8'd216;
		data_a[2721]<=8'd210;
		data_a[2722]<=8'd209;
		data_a[2723]<=8'd197;
		data_a[2724]<=8'd208;
		data_a[2725]<=8'd226;
		data_a[2726]<=8'd212;
		data_a[2727]<=8'd208;
		data_a[2728]<=8'd217;
		data_a[2729]<=8'd215;
		data_a[2730]<=8'd215;
		data_a[2731]<=8'd214;
		data_a[2732]<=8'd215;
		data_a[2733]<=8'd214;
		data_a[2734]<=8'd215;
		data_a[2735]<=8'd217;
		data_a[2736]<=8'd217;
		data_a[2737]<=8'd215;
		data_a[2738]<=8'd214;
		data_a[2739]<=8'd214;
		data_a[2740]<=8'd215;
		data_a[2741]<=8'd211;
		data_a[2742]<=8'd218;
		data_a[2743]<=8'd213;
		data_a[2744]<=8'd216;
		data_a[2745]<=8'd219;
		data_a[2746]<=8'd219;
		data_a[2747]<=8'd220;
		data_a[2748]<=8'd220;
		data_a[2749]<=8'd221;
		data_a[2750]<=8'd225;
		data_a[2751]<=8'd226;
		data_a[2752]<=8'd228;
		data_a[2753]<=8'd230;
		data_a[2754]<=8'd230;
		data_a[2755]<=8'd233;
		data_a[2756]<=8'd234;
		data_a[2757]<=8'd233;
		data_a[2758]<=8'd238;
		data_a[2759]<=8'd231;
		data_a[2760]<=8'd228;
		data_a[2761]<=8'd233;
		data_a[2762]<=8'd233;
		data_a[2763]<=8'd236;
		data_a[2764]<=8'd233;
		data_a[2765]<=8'd232;
		data_a[2766]<=8'd231;
		data_a[2767]<=8'd228;
		data_a[2768]<=8'd226;
		data_a[2769]<=8'd226;
		data_a[2770]<=8'd224;
		data_a[2771]<=8'd222;
		data_a[2772]<=8'd223;
		data_a[2773]<=8'd222;
		data_a[2774]<=8'd220;
		data_a[2775]<=8'd218;
		data_a[2776]<=8'd218;
		data_a[2777]<=8'd217;
		data_a[2778]<=8'd217;
		data_a[2779]<=8'd216;
		data_a[2780]<=8'd216;
		data_a[2781]<=8'd210;
		data_a[2782]<=8'd213;
		data_a[2783]<=8'd218;
		data_a[2784]<=8'd137;
		data_a[2785]<=8'd151;
		data_a[2786]<=8'd121;
		data_a[2787]<=8'd128;
		data_a[2788]<=8'd99;
		data_a[2789]<=8'd89;
		data_a[2790]<=8'd94;
		data_a[2791]<=8'd99;
		data_a[2792]<=8'd86;
		data_a[2793]<=8'd93;
		data_a[2794]<=8'd100;
		data_a[2795]<=8'd102;
		data_a[2796]<=8'd101;
		data_a[2797]<=8'd106;
		data_a[2798]<=8'd93;
		data_a[2799]<=8'd88;
		data_a[2800]<=8'd94;
		data_a[2801]<=8'd116;
		data_a[2802]<=8'd134;
		data_a[2803]<=8'd124;
		data_a[2804]<=8'd113;
		data_a[2805]<=8'd111;
		data_a[2806]<=8'd120;
		data_a[2807]<=8'd114;
		data_a[2808]<=8'd107;
		data_a[2809]<=8'd112;
		data_a[2810]<=8'd114;
		data_a[2811]<=8'd124;
		data_a[2812]<=8'd124;
		data_a[2813]<=8'd114;
		data_a[2814]<=8'd111;
		data_a[2815]<=8'd121;
		data_a[2816]<=8'd135;
		data_a[2817]<=8'd117;
		data_a[2818]<=8'd144;
		data_a[2819]<=8'd157;
		data_a[2820]<=8'd160;
		data_a[2821]<=8'd212;
		data_a[2822]<=8'd213;
		data_a[2823]<=8'd215;
		data_a[2824]<=8'd226;
		data_a[2825]<=8'd219;
		data_a[2826]<=8'd222;
		data_a[2827]<=8'd223;
		data_a[2828]<=8'd221;
		data_a[2829]<=8'd229;
		data_a[2830]<=8'd231;
		data_a[2831]<=8'd252;
		data_a[2832]<=8'd252;
		data_a[2833]<=8'd255;
		data_a[2834]<=8'd255;
		data_a[2835]<=8'd255;
		data_a[2836]<=8'd255;
		data_a[2837]<=8'd255;
		data_a[2838]<=8'd255;
		data_a[2839]<=8'd255;
		data_a[2840]<=8'd255;
		data_a[2841]<=8'd255;
		data_a[2842]<=8'd255;
		data_a[2843]<=8'd255;
		data_a[2844]<=8'd254;
		data_a[2845]<=8'd254;
		data_a[2846]<=8'd254;
		data_a[2847]<=8'd254;
		data_a[2848]<=8'd254;
		data_a[2849]<=8'd255;
		data_a[2850]<=8'd255;
		data_a[2851]<=8'd225;
		data_a[2852]<=8'd224;
		data_a[2853]<=8'd219;
		data_a[2854]<=8'd223;
		data_a[2855]<=8'd220;
		data_a[2856]<=8'd220;
		data_a[2857]<=8'd216;
		data_a[2858]<=8'd215;
		data_a[2859]<=8'd217;
		data_a[2860]<=8'd211;
		data_a[2861]<=8'd212;
		data_a[2862]<=8'd204;
		data_a[2863]<=8'd218;
		data_a[2864]<=8'd213;
		data_a[2865]<=8'd222;
		data_a[2866]<=8'd216;
		data_a[2867]<=8'd213;
		data_a[2868]<=8'd216;
		data_a[2869]<=8'd215;
		data_a[2870]<=8'd204;
		data_a[2871]<=8'd201;
		data_a[2872]<=8'd219;
		data_a[2873]<=8'd216;
		data_a[2874]<=8'd216;
		data_a[2875]<=8'd217;
		data_a[2876]<=8'd213;
		data_a[2877]<=8'd216;
		data_a[2878]<=8'd211;
		data_a[2879]<=8'd210;
		data_a[2880]<=8'd220;
		data_a[2881]<=8'd210;
		data_a[2882]<=8'd214;
		data_a[2883]<=8'd213;
		data_a[2884]<=8'd214;
		data_a[2885]<=8'd215;
		data_a[2886]<=8'd216;
		data_a[2887]<=8'd216;
		data_a[2888]<=8'd215;
		data_a[2889]<=8'd215;
		data_a[2890]<=8'd215;
		data_a[2891]<=8'd211;
		data_a[2892]<=8'd213;
		data_a[2893]<=8'd217;
		data_a[2894]<=8'd206;
		data_a[2895]<=8'd215;
		data_a[2896]<=8'd217;
		data_a[2897]<=8'd221;
		data_a[2898]<=8'd220;
		data_a[2899]<=8'd221;
		data_a[2900]<=8'd224;
		data_a[2901]<=8'd225;
		data_a[2902]<=8'd225;
		data_a[2903]<=8'd227;
		data_a[2904]<=8'd228;
		data_a[2905]<=8'd230;
		data_a[2906]<=8'd235;
		data_a[2907]<=8'd230;
		data_a[2908]<=8'd234;
		data_a[2909]<=8'd234;
		data_a[2910]<=8'd232;
		data_a[2911]<=8'd235;
		data_a[2912]<=8'd233;
		data_a[2913]<=8'd231;
		data_a[2914]<=8'd230;
		data_a[2915]<=8'd229;
		data_a[2916]<=8'd227;
		data_a[2917]<=8'd225;
		data_a[2918]<=8'd225;
		data_a[2919]<=8'd225;
		data_a[2920]<=8'd224;
		data_a[2921]<=8'd222;
		data_a[2922]<=8'd222;
		data_a[2923]<=8'd221;
		data_a[2924]<=8'd220;
		data_a[2925]<=8'd219;
		data_a[2926]<=8'd218;
		data_a[2927]<=8'd217;
		data_a[2928]<=8'd216;
		data_a[2929]<=8'd215;
		data_a[2930]<=8'd214;
		data_a[2931]<=8'd216;
		data_a[2932]<=8'd210;
		data_a[2933]<=8'd177;
		data_a[2934]<=8'd156;
		data_a[2935]<=8'd124;
		data_a[2936]<=8'd102;
		data_a[2937]<=8'd112;
		data_a[2938]<=8'd100;
		data_a[2939]<=8'd85;
		data_a[2940]<=8'd87;
		data_a[2941]<=8'd87;
		data_a[2942]<=8'd86;
		data_a[2943]<=8'd86;
		data_a[2944]<=8'd92;
		data_a[2945]<=8'd85;
		data_a[2946]<=8'd93;
		data_a[2947]<=8'd92;
		data_a[2948]<=8'd94;
		data_a[2949]<=8'd84;
		data_a[2950]<=8'd86;
		data_a[2951]<=8'd86;
		data_a[2952]<=8'd88;
		data_a[2953]<=8'd100;
		data_a[2954]<=8'd120;
		data_a[2955]<=8'd112;
		data_a[2956]<=8'd117;
		data_a[2957]<=8'd111;
		data_a[2958]<=8'd108;
		data_a[2959]<=8'd110;
		data_a[2960]<=8'd105;
		data_a[2961]<=8'd111;
		data_a[2962]<=8'd120;
		data_a[2963]<=8'd115;
		data_a[2964]<=8'd110;
		data_a[2965]<=8'd111;
		data_a[2966]<=8'd129;
		data_a[2967]<=8'd124;
		data_a[2968]<=8'd138;
		data_a[2969]<=8'd158;
		data_a[2970]<=8'd159;
		data_a[2971]<=8'd174;
		data_a[2972]<=8'd216;
		data_a[2973]<=8'd223;
		data_a[2974]<=8'd218;
		data_a[2975]<=8'd216;
		data_a[2976]<=8'd223;
		data_a[2977]<=8'd222;
		data_a[2978]<=8'd223;
		data_a[2979]<=8'd229;
		data_a[2980]<=8'd230;
		data_a[2981]<=8'd244;
		data_a[2982]<=8'd253;
		data_a[2983]<=8'd255;
		data_a[2984]<=8'd255;
		data_a[2985]<=8'd255;
		data_a[2986]<=8'd255;
		data_a[2987]<=8'd255;
		data_a[2988]<=8'd255;
		data_a[2989]<=8'd255;
		data_a[2990]<=8'd255;
		data_a[2991]<=8'd255;
		data_a[2992]<=8'd255;
		data_a[2993]<=8'd255;
		data_a[2994]<=8'd254;
		data_a[2995]<=8'd254;
		data_a[2996]<=8'd254;
		data_a[2997]<=8'd254;
		data_a[2998]<=8'd254;
		data_a[2999]<=8'd254;
		data_a[3000]<=8'd254;
		data_a[3001]<=8'd224;
		data_a[3002]<=8'd222;
		data_a[3003]<=8'd223;
		data_a[3004]<=8'd222;
		data_a[3005]<=8'd220;
		data_a[3006]<=8'd216;
		data_a[3007]<=8'd216;
		data_a[3008]<=8'd216;
		data_a[3009]<=8'd213;
		data_a[3010]<=8'd216;
		data_a[3011]<=8'd221;
		data_a[3012]<=8'd208;
		data_a[3013]<=8'd198;
		data_a[3014]<=8'd219;
		data_a[3015]<=8'd213;
		data_a[3016]<=8'd219;
		data_a[3017]<=8'd219;
		data_a[3018]<=8'd205;
		data_a[3019]<=8'd201;
		data_a[3020]<=8'd215;
		data_a[3021]<=8'd212;
		data_a[3022]<=8'd211;
		data_a[3023]<=8'd213;
		data_a[3024]<=8'd214;
		data_a[3025]<=8'd207;
		data_a[3026]<=8'd210;
		data_a[3027]<=8'd217;
		data_a[3028]<=8'd215;
		data_a[3029]<=8'd210;
		data_a[3030]<=8'd213;
		data_a[3031]<=8'd213;
		data_a[3032]<=8'd214;
		data_a[3033]<=8'd212;
		data_a[3034]<=8'd212;
		data_a[3035]<=8'd213;
		data_a[3036]<=8'd215;
		data_a[3037]<=8'd215;
		data_a[3038]<=8'd215;
		data_a[3039]<=8'd215;
		data_a[3040]<=8'd215;
		data_a[3041]<=8'd219;
		data_a[3042]<=8'd210;
		data_a[3043]<=8'd217;
		data_a[3044]<=8'd213;
		data_a[3045]<=8'd217;
		data_a[3046]<=8'd217;
		data_a[3047]<=8'd222;
		data_a[3048]<=8'd220;
		data_a[3049]<=8'd222;
		data_a[3050]<=8'd222;
		data_a[3051]<=8'd224;
		data_a[3052]<=8'd225;
		data_a[3053]<=8'd226;
		data_a[3054]<=8'd228;
		data_a[3055]<=8'd229;
		data_a[3056]<=8'd232;
		data_a[3057]<=8'd232;
		data_a[3058]<=8'd233;
		data_a[3059]<=8'd236;
		data_a[3060]<=8'd230;
		data_a[3061]<=8'd225;
		data_a[3062]<=8'd231;
		data_a[3063]<=8'd231;
		data_a[3064]<=8'd229;
		data_a[3065]<=8'd228;
		data_a[3066]<=8'd226;
		data_a[3067]<=8'd224;
		data_a[3068]<=8'd224;
		data_a[3069]<=8'd225;
		data_a[3070]<=8'd224;
		data_a[3071]<=8'd222;
		data_a[3072]<=8'd220;
		data_a[3073]<=8'd219;
		data_a[3074]<=8'd218;
		data_a[3075]<=8'd217;
		data_a[3076]<=8'd216;
		data_a[3077]<=8'd216;
		data_a[3078]<=8'd215;
		data_a[3079]<=8'd215;
		data_a[3080]<=8'd217;
		data_a[3081]<=8'd209;
		data_a[3082]<=8'd158;
		data_a[3083]<=8'd137;
		data_a[3084]<=8'd104;
		data_a[3085]<=8'd108;
		data_a[3086]<=8'd97;
		data_a[3087]<=8'd100;
		data_a[3088]<=8'd104;
		data_a[3089]<=8'd94;
		data_a[3090]<=8'd87;
		data_a[3091]<=8'd82;
		data_a[3092]<=8'd83;
		data_a[3093]<=8'd80;
		data_a[3094]<=8'd84;
		data_a[3095]<=8'd80;
		data_a[3096]<=8'd78;
		data_a[3097]<=8'd81;
		data_a[3098]<=8'd92;
		data_a[3099]<=8'd87;
		data_a[3100]<=8'd79;
		data_a[3101]<=8'd75;
		data_a[3102]<=8'd85;
		data_a[3103]<=8'd86;
		data_a[3104]<=8'd91;
		data_a[3105]<=8'd99;
		data_a[3106]<=8'd107;
		data_a[3107]<=8'd110;
		data_a[3108]<=8'd116;
		data_a[3109]<=8'd119;
		data_a[3110]<=8'd112;
		data_a[3111]<=8'd104;
		data_a[3112]<=8'd108;
		data_a[3113]<=8'd113;
		data_a[3114]<=8'd112;
		data_a[3115]<=8'd107;
		data_a[3116]<=8'd129;
		data_a[3117]<=8'd126;
		data_a[3118]<=8'd129;
		data_a[3119]<=8'd154;
		data_a[3120]<=8'd158;
		data_a[3121]<=8'd149;
		data_a[3122]<=8'd187;
		data_a[3123]<=8'd219;
		data_a[3124]<=8'd222;
		data_a[3125]<=8'd218;
		data_a[3126]<=8'd219;
		data_a[3127]<=8'd228;
		data_a[3128]<=8'd225;
		data_a[3129]<=8'd225;
		data_a[3130]<=8'd228;
		data_a[3131]<=8'd237;
		data_a[3132]<=8'd255;
		data_a[3133]<=8'd254;
		data_a[3134]<=8'd255;
		data_a[3135]<=8'd255;
		data_a[3136]<=8'd255;
		data_a[3137]<=8'd255;
		data_a[3138]<=8'd255;
		data_a[3139]<=8'd255;
		data_a[3140]<=8'd255;
		data_a[3141]<=8'd255;
		data_a[3142]<=8'd255;
		data_a[3143]<=8'd255;
		data_a[3144]<=8'd255;
		data_a[3145]<=8'd255;
		data_a[3146]<=8'd254;
		data_a[3147]<=8'd254;
		data_a[3148]<=8'd255;
		data_a[3149]<=8'd255;
		data_a[3150]<=8'd254;
		data_a[3151]<=8'd219;
		data_a[3152]<=8'd225;
		data_a[3153]<=8'd223;
		data_a[3154]<=8'd217;
		data_a[3155]<=8'd221;
		data_a[3156]<=8'd215;
		data_a[3157]<=8'd222;
		data_a[3158]<=8'd214;
		data_a[3159]<=8'd216;
		data_a[3160]<=8'd217;
		data_a[3161]<=8'd212;
		data_a[3162]<=8'd213;
		data_a[3163]<=8'd220;
		data_a[3164]<=8'd193;
		data_a[3165]<=8'd206;
		data_a[3166]<=8'd200;
		data_a[3167]<=8'd206;
		data_a[3168]<=8'd214;
		data_a[3169]<=8'd211;
		data_a[3170]<=8'd213;
		data_a[3171]<=8'd213;
		data_a[3172]<=8'd216;
		data_a[3173]<=8'd214;
		data_a[3174]<=8'd217;
		data_a[3175]<=8'd215;
		data_a[3176]<=8'd217;
		data_a[3177]<=8'd212;
		data_a[3178]<=8'd211;
		data_a[3179]<=8'd216;
		data_a[3180]<=8'd213;
		data_a[3181]<=8'd211;
		data_a[3182]<=8'd215;
		data_a[3183]<=8'd213;
		data_a[3184]<=8'd212;
		data_a[3185]<=8'd213;
		data_a[3186]<=8'd215;
		data_a[3187]<=8'd215;
		data_a[3188]<=8'd215;
		data_a[3189]<=8'd214;
		data_a[3190]<=8'd211;
		data_a[3191]<=8'd210;
		data_a[3192]<=8'd205;
		data_a[3193]<=8'd211;
		data_a[3194]<=8'd212;
		data_a[3195]<=8'd215;
		data_a[3196]<=8'd221;
		data_a[3197]<=8'd213;
		data_a[3198]<=8'd220;
		data_a[3199]<=8'd221;
		data_a[3200]<=8'd220;
		data_a[3201]<=8'd223;
		data_a[3202]<=8'd225;
		data_a[3203]<=8'd226;
		data_a[3204]<=8'd229;
		data_a[3205]<=8'd228;
		data_a[3206]<=8'd229;
		data_a[3207]<=8'd232;
		data_a[3208]<=8'd229;
		data_a[3209]<=8'd231;
		data_a[3210]<=8'd225;
		data_a[3211]<=8'd219;
		data_a[3212]<=8'd228;
		data_a[3213]<=8'd231;
		data_a[3214]<=8'd228;
		data_a[3215]<=8'd228;
		data_a[3216]<=8'd227;
		data_a[3217]<=8'd225;
		data_a[3218]<=8'd224;
		data_a[3219]<=8'd224;
		data_a[3220]<=8'd223;
		data_a[3221]<=8'd222;
		data_a[3222]<=8'd219;
		data_a[3223]<=8'd218;
		data_a[3224]<=8'd217;
		data_a[3225]<=8'd216;
		data_a[3226]<=8'd215;
		data_a[3227]<=8'd215;
		data_a[3228]<=8'd216;
		data_a[3229]<=8'd216;
		data_a[3230]<=8'd212;
		data_a[3231]<=8'd171;
		data_a[3232]<=8'd123;
		data_a[3233]<=8'd116;
		data_a[3234]<=8'd112;
		data_a[3235]<=8'd108;
		data_a[3236]<=8'd96;
		data_a[3237]<=8'd89;
		data_a[3238]<=8'd83;
		data_a[3239]<=8'd92;
		data_a[3240]<=8'd87;
		data_a[3241]<=8'd87;
		data_a[3242]<=8'd82;
		data_a[3243]<=8'd80;
		data_a[3244]<=8'd77;
		data_a[3245]<=8'd80;
		data_a[3246]<=8'd77;
		data_a[3247]<=8'd80;
		data_a[3248]<=8'd70;
		data_a[3249]<=8'd77;
		data_a[3250]<=8'd81;
		data_a[3251]<=8'd71;
		data_a[3252]<=8'd86;
		data_a[3253]<=8'd78;
		data_a[3254]<=8'd79;
		data_a[3255]<=8'd87;
		data_a[3256]<=8'd87;
		data_a[3257]<=8'd92;
		data_a[3258]<=8'd97;
		data_a[3259]<=8'd99;
		data_a[3260]<=8'd103;
		data_a[3261]<=8'd102;
		data_a[3262]<=8'd98;
		data_a[3263]<=8'd106;
		data_a[3264]<=8'd110;
		data_a[3265]<=8'd111;
		data_a[3266]<=8'd132;
		data_a[3267]<=8'd110;
		data_a[3268]<=8'd119;
		data_a[3269]<=8'd142;
		data_a[3270]<=8'd161;
		data_a[3271]<=8'd141;
		data_a[3272]<=8'd157;
		data_a[3273]<=8'd219;
		data_a[3274]<=8'd220;
		data_a[3275]<=8'd218;
		data_a[3276]<=8'd228;
		data_a[3277]<=8'd222;
		data_a[3278]<=8'd225;
		data_a[3279]<=8'd224;
		data_a[3280]<=8'd228;
		data_a[3281]<=8'd235;
		data_a[3282]<=8'd254;
		data_a[3283]<=8'd254;
		data_a[3284]<=8'd255;
		data_a[3285]<=8'd255;
		data_a[3286]<=8'd255;
		data_a[3287]<=8'd255;
		data_a[3288]<=8'd255;
		data_a[3289]<=8'd255;
		data_a[3290]<=8'd255;
		data_a[3291]<=8'd255;
		data_a[3292]<=8'd255;
		data_a[3293]<=8'd255;
		data_a[3294]<=8'd255;
		data_a[3295]<=8'd254;
		data_a[3296]<=8'd254;
		data_a[3297]<=8'd254;
		data_a[3298]<=8'd255;
		data_a[3299]<=8'd255;
		data_a[3300]<=8'd254;
		data_a[3301]<=8'd176;
		data_a[3302]<=8'd213;
		data_a[3303]<=8'd222;
		data_a[3304]<=8'd213;
		data_a[3305]<=8'd218;
		data_a[3306]<=8'd215;
		data_a[3307]<=8'd213;
		data_a[3308]<=8'd217;
		data_a[3309]<=8'd213;
		data_a[3310]<=8'd212;
		data_a[3311]<=8'd215;
		data_a[3312]<=8'd214;
		data_a[3313]<=8'd212;
		data_a[3314]<=8'd224;
		data_a[3315]<=8'd194;
		data_a[3316]<=8'd213;
		data_a[3317]<=8'd214;
		data_a[3318]<=8'd217;
		data_a[3319]<=8'd210;
		data_a[3320]<=8'd215;
		data_a[3321]<=8'd216;
		data_a[3322]<=8'd211;
		data_a[3323]<=8'd215;
		data_a[3324]<=8'd213;
		data_a[3325]<=8'd211;
		data_a[3326]<=8'd214;
		data_a[3327]<=8'd215;
		data_a[3328]<=8'd216;
		data_a[3329]<=8'd214;
		data_a[3330]<=8'd209;
		data_a[3331]<=8'd211;
		data_a[3332]<=8'd214;
		data_a[3333]<=8'd212;
		data_a[3334]<=8'd211;
		data_a[3335]<=8'd212;
		data_a[3336]<=8'd214;
		data_a[3337]<=8'd213;
		data_a[3338]<=8'd212;
		data_a[3339]<=8'd211;
		data_a[3340]<=8'd202;
		data_a[3341]<=8'd223;
		data_a[3342]<=8'd204;
		data_a[3343]<=8'd193;
		data_a[3344]<=8'd214;
		data_a[3345]<=8'd220;
		data_a[3346]<=8'd210;
		data_a[3347]<=8'd221;
		data_a[3348]<=8'd217;
		data_a[3349]<=8'd219;
		data_a[3350]<=8'd217;
		data_a[3351]<=8'd222;
		data_a[3352]<=8'd224;
		data_a[3353]<=8'd224;
		data_a[3354]<=8'd226;
		data_a[3355]<=8'd223;
		data_a[3356]<=8'd228;
		data_a[3357]<=8'd227;
		data_a[3358]<=8'd222;
		data_a[3359]<=8'd223;
		data_a[3360]<=8'd228;
		data_a[3361]<=8'd230;
		data_a[3362]<=8'd228;
		data_a[3363]<=8'd224;
		data_a[3364]<=8'd226;
		data_a[3365]<=8'd227;
		data_a[3366]<=8'd227;
		data_a[3367]<=8'd225;
		data_a[3368]<=8'd224;
		data_a[3369]<=8'd223;
		data_a[3370]<=8'd223;
		data_a[3371]<=8'd221;
		data_a[3372]<=8'd220;
		data_a[3373]<=8'd219;
		data_a[3374]<=8'd218;
		data_a[3375]<=8'd217;
		data_a[3376]<=8'd217;
		data_a[3377]<=8'd216;
		data_a[3378]<=8'd214;
		data_a[3379]<=8'd212;
		data_a[3380]<=8'd200;
		data_a[3381]<=8'd137;
		data_a[3382]<=8'd117;
		data_a[3383]<=8'd118;
		data_a[3384]<=8'd112;
		data_a[3385]<=8'd121;
		data_a[3386]<=8'd124;
		data_a[3387]<=8'd89;
		data_a[3388]<=8'd77;
		data_a[3389]<=8'd86;
		data_a[3390]<=8'd79;
		data_a[3391]<=8'd80;
		data_a[3392]<=8'd81;
		data_a[3393]<=8'd84;
		data_a[3394]<=8'd80;
		data_a[3395]<=8'd76;
		data_a[3396]<=8'd72;
		data_a[3397]<=8'd75;
		data_a[3398]<=8'd78;
		data_a[3399]<=8'd73;
		data_a[3400]<=8'd78;
		data_a[3401]<=8'd78;
		data_a[3402]<=8'd74;
		data_a[3403]<=8'd75;
		data_a[3404]<=8'd80;
		data_a[3405]<=8'd82;
		data_a[3406]<=8'd80;
		data_a[3407]<=8'd85;
		data_a[3408]<=8'd89;
		data_a[3409]<=8'd86;
		data_a[3410]<=8'd94;
		data_a[3411]<=8'd104;
		data_a[3412]<=8'd100;
		data_a[3413]<=8'd98;
		data_a[3414]<=8'd100;
		data_a[3415]<=8'd110;
		data_a[3416]<=8'd126;
		data_a[3417]<=8'd108;
		data_a[3418]<=8'd115;
		data_a[3419]<=8'd125;
		data_a[3420]<=8'd139;
		data_a[3421]<=8'd139;
		data_a[3422]<=8'd176;
		data_a[3423]<=8'd212;
		data_a[3424]<=8'd219;
		data_a[3425]<=8'd223;
		data_a[3426]<=8'd214;
		data_a[3427]<=8'd227;
		data_a[3428]<=8'd223;
		data_a[3429]<=8'd225;
		data_a[3430]<=8'd228;
		data_a[3431]<=8'd234;
		data_a[3432]<=8'd246;
		data_a[3433]<=8'd255;
		data_a[3434]<=8'd255;
		data_a[3435]<=8'd255;
		data_a[3436]<=8'd255;
		data_a[3437]<=8'd255;
		data_a[3438]<=8'd255;
		data_a[3439]<=8'd255;
		data_a[3440]<=8'd255;
		data_a[3441]<=8'd255;
		data_a[3442]<=8'd255;
		data_a[3443]<=8'd255;
		data_a[3444]<=8'd255;
		data_a[3445]<=8'd255;
		data_a[3446]<=8'd255;
		data_a[3447]<=8'd254;
		data_a[3448]<=8'd253;
		data_a[3449]<=8'd252;
		data_a[3450]<=8'd254;
		data_a[3451]<=8'd190;
		data_a[3452]<=8'd121;
		data_a[3453]<=8'd208;
		data_a[3454]<=8'd220;
		data_a[3455]<=8'd215;
		data_a[3456]<=8'd215;
		data_a[3457]<=8'd217;
		data_a[3458]<=8'd215;
		data_a[3459]<=8'd214;
		data_a[3460]<=8'd218;
		data_a[3461]<=8'd212;
		data_a[3462]<=8'd215;
		data_a[3463]<=8'd217;
		data_a[3464]<=8'd217;
		data_a[3465]<=8'd223;
		data_a[3466]<=8'd216;
		data_a[3467]<=8'd203;
		data_a[3468]<=8'd215;
		data_a[3469]<=8'd214;
		data_a[3470]<=8'd214;
		data_a[3471]<=8'd215;
		data_a[3472]<=8'd213;
		data_a[3473]<=8'd216;
		data_a[3474]<=8'd214;
		data_a[3475]<=8'd211;
		data_a[3476]<=8'd213;
		data_a[3477]<=8'd215;
		data_a[3478]<=8'd212;
		data_a[3479]<=8'd210;
		data_a[3480]<=8'd212;
		data_a[3481]<=8'd210;
		data_a[3482]<=8'd211;
		data_a[3483]<=8'd209;
		data_a[3484]<=8'd208;
		data_a[3485]<=8'd209;
		data_a[3486]<=8'd211;
		data_a[3487]<=8'd209;
		data_a[3488]<=8'd207;
		data_a[3489]<=8'd205;
		data_a[3490]<=8'd200;
		data_a[3491]<=8'd195;
		data_a[3492]<=8'd196;
		data_a[3493]<=8'd191;
		data_a[3494]<=8'd170;
		data_a[3495]<=8'd204;
		data_a[3496]<=8'd214;
		data_a[3497]<=8'd204;
		data_a[3498]<=8'd214;
		data_a[3499]<=8'd217;
		data_a[3500]<=8'd214;
		data_a[3501]<=8'd220;
		data_a[3502]<=8'd223;
		data_a[3503]<=8'd221;
		data_a[3504]<=8'd222;
		data_a[3505]<=8'd217;
		data_a[3506]<=8'd214;
		data_a[3507]<=8'd223;
		data_a[3508]<=8'd231;
		data_a[3509]<=8'd225;
		data_a[3510]<=8'd228;
		data_a[3511]<=8'd232;
		data_a[3512]<=8'd227;
		data_a[3513]<=8'd229;
		data_a[3514]<=8'd223;
		data_a[3515]<=8'd225;
		data_a[3516]<=8'd226;
		data_a[3517]<=8'd225;
		data_a[3518]<=8'd224;
		data_a[3519]<=8'd223;
		data_a[3520]<=8'd222;
		data_a[3521]<=8'd222;
		data_a[3522]<=8'd220;
		data_a[3523]<=8'd219;
		data_a[3524]<=8'd218;
		data_a[3525]<=8'd219;
		data_a[3526]<=8'd218;
		data_a[3527]<=8'd215;
		data_a[3528]<=8'd210;
		data_a[3529]<=8'd205;
		data_a[3530]<=8'd131;
		data_a[3531]<=8'd137;
		data_a[3532]<=8'd128;
		data_a[3533]<=8'd113;
		data_a[3534]<=8'd124;
		data_a[3535]<=8'd111;
		data_a[3536]<=8'd107;
		data_a[3537]<=8'd106;
		data_a[3538]<=8'd99;
		data_a[3539]<=8'd103;
		data_a[3540]<=8'd98;
		data_a[3541]<=8'd87;
		data_a[3542]<=8'd84;
		data_a[3543]<=8'd78;
		data_a[3544]<=8'd78;
		data_a[3545]<=8'd67;
		data_a[3546]<=8'd73;
		data_a[3547]<=8'd71;
		data_a[3548]<=8'd74;
		data_a[3549]<=8'd78;
		data_a[3550]<=8'd73;
		data_a[3551]<=8'd73;
		data_a[3552]<=8'd81;
		data_a[3553]<=8'd76;
		data_a[3554]<=8'd77;
		data_a[3555]<=8'd82;
		data_a[3556]<=8'd83;
		data_a[3557]<=8'd82;
		data_a[3558]<=8'd85;
		data_a[3559]<=8'd87;
		data_a[3560]<=8'd88;
		data_a[3561]<=8'd95;
		data_a[3562]<=8'd98;
		data_a[3563]<=8'd96;
		data_a[3564]<=8'd101;
		data_a[3565]<=8'd109;
		data_a[3566]<=8'd109;
		data_a[3567]<=8'd111;
		data_a[3568]<=8'd116;
		data_a[3569]<=8'd124;
		data_a[3570]<=8'd142;
		data_a[3571]<=8'd150;
		data_a[3572]<=8'd201;
		data_a[3573]<=8'd212;
		data_a[3574]<=8'd216;
		data_a[3575]<=8'd221;
		data_a[3576]<=8'd223;
		data_a[3577]<=8'd223;
		data_a[3578]<=8'd221;
		data_a[3579]<=8'd227;
		data_a[3580]<=8'd227;
		data_a[3581]<=8'd234;
		data_a[3582]<=8'd237;
		data_a[3583]<=8'd254;
		data_a[3584]<=8'd254;
		data_a[3585]<=8'd255;
		data_a[3586]<=8'd255;
		data_a[3587]<=8'd255;
		data_a[3588]<=8'd255;
		data_a[3589]<=8'd255;
		data_a[3590]<=8'd255;
		data_a[3591]<=8'd255;
		data_a[3592]<=8'd255;
		data_a[3593]<=8'd255;
		data_a[3594]<=8'd252;
		data_a[3595]<=8'd253;
		data_a[3596]<=8'd251;
		data_a[3597]<=8'd247;
		data_a[3598]<=8'd241;
		data_a[3599]<=8'd237;
		data_a[3600]<=8'd254;
		data_a[3601]<=8'd205;
		data_a[3602]<=8'd193;
		data_a[3603]<=8'd100;
		data_a[3604]<=8'd189;
		data_a[3605]<=8'd220;
		data_a[3606]<=8'd215;
		data_a[3607]<=8'd219;
		data_a[3608]<=8'd213;
		data_a[3609]<=8'd216;
		data_a[3610]<=8'd217;
		data_a[3611]<=8'd209;
		data_a[3612]<=8'd218;
		data_a[3613]<=8'd213;
		data_a[3614]<=8'd211;
		data_a[3615]<=8'd218;
		data_a[3616]<=8'd212;
		data_a[3617]<=8'd213;
		data_a[3618]<=8'd204;
		data_a[3619]<=8'd216;
		data_a[3620]<=8'd215;
		data_a[3621]<=8'd217;
		data_a[3622]<=8'd211;
		data_a[3623]<=8'd212;
		data_a[3624]<=8'd212;
		data_a[3625]<=8'd213;
		data_a[3626]<=8'd216;
		data_a[3627]<=8'd206;
		data_a[3628]<=8'd213;
		data_a[3629]<=8'd210;
		data_a[3630]<=8'd213;
		data_a[3631]<=8'd210;
		data_a[3632]<=8'd213;
		data_a[3633]<=8'd207;
		data_a[3634]<=8'd211;
		data_a[3635]<=8'd211;
		data_a[3636]<=8'd219;
		data_a[3637]<=8'd188;
		data_a[3638]<=8'd189;
		data_a[3639]<=8'd197;
		data_a[3640]<=8'd158;
		data_a[3641]<=8'd136;
		data_a[3642]<=8'd165;
		data_a[3643]<=8'd156;
		data_a[3644]<=8'd142;
		data_a[3645]<=8'd182;
		data_a[3646]<=8'd187;
		data_a[3647]<=8'd211;
		data_a[3648]<=8'd213;
		data_a[3649]<=8'd200;
		data_a[3650]<=8'd219;
		data_a[3651]<=8'd210;
		data_a[3652]<=8'd220;
		data_a[3653]<=8'd209;
		data_a[3654]<=8'd209;
		data_a[3655]<=8'd222;
		data_a[3656]<=8'd225;
		data_a[3657]<=8'd226;
		data_a[3658]<=8'd222;
		data_a[3659]<=8'd225;
		data_a[3660]<=8'd225;
		data_a[3661]<=8'd228;
		data_a[3662]<=8'd225;
		data_a[3663]<=8'd230;
		data_a[3664]<=8'd223;
		data_a[3665]<=8'd220;
		data_a[3666]<=8'd221;
		data_a[3667]<=8'd224;
		data_a[3668]<=8'd225;
		data_a[3669]<=8'd220;
		data_a[3670]<=8'd227;
		data_a[3671]<=8'd219;
		data_a[3672]<=8'd219;
		data_a[3673]<=8'd217;
		data_a[3674]<=8'd214;
		data_a[3675]<=8'd209;
		data_a[3676]<=8'd208;
		data_a[3677]<=8'd214;
		data_a[3678]<=8'd211;
		data_a[3679]<=8'd158;
		data_a[3680]<=8'd129;
		data_a[3681]<=8'd141;
		data_a[3682]<=8'd113;
		data_a[3683]<=8'd115;
		data_a[3684]<=8'd103;
		data_a[3685]<=8'd115;
		data_a[3686]<=8'd115;
		data_a[3687]<=8'd117;
		data_a[3688]<=8'd115;
		data_a[3689]<=8'd105;
		data_a[3690]<=8'd94;
		data_a[3691]<=8'd95;
		data_a[3692]<=8'd90;
		data_a[3693]<=8'd86;
		data_a[3694]<=8'd77;
		data_a[3695]<=8'd74;
		data_a[3696]<=8'd70;
		data_a[3697]<=8'd73;
		data_a[3698]<=8'd71;
		data_a[3699]<=8'd70;
		data_a[3700]<=8'd75;
		data_a[3701]<=8'd73;
		data_a[3702]<=8'd75;
		data_a[3703]<=8'd73;
		data_a[3704]<=8'd73;
		data_a[3705]<=8'd78;
		data_a[3706]<=8'd82;
		data_a[3707]<=8'd86;
		data_a[3708]<=8'd90;
		data_a[3709]<=8'd90;
		data_a[3710]<=8'd88;
		data_a[3711]<=8'd89;
		data_a[3712]<=8'd96;
		data_a[3713]<=8'd89;
		data_a[3714]<=8'd103;
		data_a[3715]<=8'd106;
		data_a[3716]<=8'd104;
		data_a[3717]<=8'd107;
		data_a[3718]<=8'd117;
		data_a[3719]<=8'd119;
		data_a[3720]<=8'd134;
		data_a[3721]<=8'd145;
		data_a[3722]<=8'd192;
		data_a[3723]<=8'd189;
		data_a[3724]<=8'd196;
		data_a[3725]<=8'd223;
		data_a[3726]<=8'd219;
		data_a[3727]<=8'd220;
		data_a[3728]<=8'd224;
		data_a[3729]<=8'd223;
		data_a[3730]<=8'd226;
		data_a[3731]<=8'd234;
		data_a[3732]<=8'd238;
		data_a[3733]<=8'd251;
		data_a[3734]<=8'd253;
		data_a[3735]<=8'd254;
		data_a[3736]<=8'd254;
		data_a[3737]<=8'd254;
		data_a[3738]<=8'd254;
		data_a[3739]<=8'd254;
		data_a[3740]<=8'd254;
		data_a[3741]<=8'd253;
		data_a[3742]<=8'd252;
		data_a[3743]<=8'd248;
		data_a[3744]<=8'd245;
		data_a[3745]<=8'd243;
		data_a[3746]<=8'd240;
		data_a[3747]<=8'd238;
		data_a[3748]<=8'd236;
		data_a[3749]<=8'd235;
		data_a[3750]<=8'd254;
		data_a[3751]<=8'd122;
		data_a[3752]<=8'd229;
		data_a[3753]<=8'd198;
		data_a[3754]<=8'd115;
		data_a[3755]<=8'd149;
		data_a[3756]<=8'd203;
		data_a[3757]<=8'd225;
		data_a[3758]<=8'd213;
		data_a[3759]<=8'd211;
		data_a[3760]<=8'd216;
		data_a[3761]<=8'd215;
		data_a[3762]<=8'd214;
		data_a[3763]<=8'd213;
		data_a[3764]<=8'd216;
		data_a[3765]<=8'd211;
		data_a[3766]<=8'd212;
		data_a[3767]<=8'd208;
		data_a[3768]<=8'd212;
		data_a[3769]<=8'd198;
		data_a[3770]<=8'd217;
		data_a[3771]<=8'd215;
		data_a[3772]<=8'd215;
		data_a[3773]<=8'd212;
		data_a[3774]<=8'd212;
		data_a[3775]<=8'd211;
		data_a[3776]<=8'd212;
		data_a[3777]<=8'd213;
		data_a[3778]<=8'd213;
		data_a[3779]<=8'd211;
		data_a[3780]<=8'd209;
		data_a[3781]<=8'd208;
		data_a[3782]<=8'd213;
		data_a[3783]<=8'd210;
		data_a[3784]<=8'd182;
		data_a[3785]<=8'd184;
		data_a[3786]<=8'd128;
		data_a[3787]<=8'd125;
		data_a[3788]<=8'd152;
		data_a[3789]<=8'd163;
		data_a[3790]<=8'd179;
		data_a[3791]<=8'd193;
		data_a[3792]<=8'd128;
		data_a[3793]<=8'd114;
		data_a[3794]<=8'd107;
		data_a[3795]<=8'd126;
		data_a[3796]<=8'd190;
		data_a[3797]<=8'd182;
		data_a[3798]<=8'd190;
		data_a[3799]<=8'd142;
		data_a[3800]<=8'd162;
		data_a[3801]<=8'd179;
		data_a[3802]<=8'd207;
		data_a[3803]<=8'd209;
		data_a[3804]<=8'd188;
		data_a[3805]<=8'd210;
		data_a[3806]<=8'd211;
		data_a[3807]<=8'd228;
		data_a[3808]<=8'd225;
		data_a[3809]<=8'd225;
		data_a[3810]<=8'd225;
		data_a[3811]<=8'd223;
		data_a[3812]<=8'd224;
		data_a[3813]<=8'd220;
		data_a[3814]<=8'd223;
		data_a[3815]<=8'd225;
		data_a[3816]<=8'd225;
		data_a[3817]<=8'd223;
		data_a[3818]<=8'd220;
		data_a[3819]<=8'd220;
		data_a[3820]<=8'd219;
		data_a[3821]<=8'd222;
		data_a[3822]<=8'd214;
		data_a[3823]<=8'd211;
		data_a[3824]<=8'd208;
		data_a[3825]<=8'd219;
		data_a[3826]<=8'd211;
		data_a[3827]<=8'd212;
		data_a[3828]<=8'd210;
		data_a[3829]<=8'd152;
		data_a[3830]<=8'd126;
		data_a[3831]<=8'd117;
		data_a[3832]<=8'd117;
		data_a[3833]<=8'd108;
		data_a[3834]<=8'd105;
		data_a[3835]<=8'd113;
		data_a[3836]<=8'd106;
		data_a[3837]<=8'd101;
		data_a[3838]<=8'd100;
		data_a[3839]<=8'd109;
		data_a[3840]<=8'd110;
		data_a[3841]<=8'd95;
		data_a[3842]<=8'd79;
		data_a[3843]<=8'd71;
		data_a[3844]<=8'd72;
		data_a[3845]<=8'd74;
		data_a[3846]<=8'd70;
		data_a[3847]<=8'd72;
		data_a[3848]<=8'd72;
		data_a[3849]<=8'd71;
		data_a[3850]<=8'd78;
		data_a[3851]<=8'd76;
		data_a[3852]<=8'd79;
		data_a[3853]<=8'd77;
		data_a[3854]<=8'd83;
		data_a[3855]<=8'd84;
		data_a[3856]<=8'd83;
		data_a[3857]<=8'd82;
		data_a[3858]<=8'd85;
		data_a[3859]<=8'd87;
		data_a[3860]<=8'd89;
		data_a[3861]<=8'd93;
		data_a[3862]<=8'd99;
		data_a[3863]<=8'd94;
		data_a[3864]<=8'd96;
		data_a[3865]<=8'd96;
		data_a[3866]<=8'd95;
		data_a[3867]<=8'd103;
		data_a[3868]<=8'd111;
		data_a[3869]<=8'd121;
		data_a[3870]<=8'd125;
		data_a[3871]<=8'd148;
		data_a[3872]<=8'd173;
		data_a[3873]<=8'd155;
		data_a[3874]<=8'd200;
		data_a[3875]<=8'd221;
		data_a[3876]<=8'd219;
		data_a[3877]<=8'd221;
		data_a[3878]<=8'd225;
		data_a[3879]<=8'd228;
		data_a[3880]<=8'd227;
		data_a[3881]<=8'd232;
		data_a[3882]<=8'd232;
		data_a[3883]<=8'd239;
		data_a[3884]<=8'd252;
		data_a[3885]<=8'd254;
		data_a[3886]<=8'd254;
		data_a[3887]<=8'd254;
		data_a[3888]<=8'd254;
		data_a[3889]<=8'd252;
		data_a[3890]<=8'd247;
		data_a[3891]<=8'd244;
		data_a[3892]<=8'd241;
		data_a[3893]<=8'd241;
		data_a[3894]<=8'd242;
		data_a[3895]<=8'd241;
		data_a[3896]<=8'd238;
		data_a[3897]<=8'd236;
		data_a[3898]<=8'd234;
		data_a[3899]<=8'd232;
		data_a[3900]<=8'd254;
		data_a[3901]<=8'd214;
		data_a[3902]<=8'd185;
		data_a[3903]<=8'd197;
		data_a[3904]<=8'd152;
		data_a[3905]<=8'd122;
		data_a[3906]<=8'd106;
		data_a[3907]<=8'd196;
		data_a[3908]<=8'd212;
		data_a[3909]<=8'd212;
		data_a[3910]<=8'd215;
		data_a[3911]<=8'd216;
		data_a[3912]<=8'd210;
		data_a[3913]<=8'd211;
		data_a[3914]<=8'd218;
		data_a[3915]<=8'd216;
		data_a[3916]<=8'd211;
		data_a[3917]<=8'd215;
		data_a[3918]<=8'd213;
		data_a[3919]<=8'd207;
		data_a[3920]<=8'd194;
		data_a[3921]<=8'd211;
		data_a[3922]<=8'd209;
		data_a[3923]<=8'd209;
		data_a[3924]<=8'd209;
		data_a[3925]<=8'd210;
		data_a[3926]<=8'd209;
		data_a[3927]<=8'd210;
		data_a[3928]<=8'd208;
		data_a[3929]<=8'd212;
		data_a[3930]<=8'd209;
		data_a[3931]<=8'd204;
		data_a[3932]<=8'd206;
		data_a[3933]<=8'd188;
		data_a[3934]<=8'd178;
		data_a[3935]<=8'd142;
		data_a[3936]<=8'd148;
		data_a[3937]<=8'd145;
		data_a[3938]<=8'd140;
		data_a[3939]<=8'd158;
		data_a[3940]<=8'd153;
		data_a[3941]<=8'd157;
		data_a[3942]<=8'd134;
		data_a[3943]<=8'd124;
		data_a[3944]<=8'd116;
		data_a[3945]<=8'd101;
		data_a[3946]<=8'd134;
		data_a[3947]<=8'd163;
		data_a[3948]<=8'd142;
		data_a[3949]<=8'd172;
		data_a[3950]<=8'd175;
		data_a[3951]<=8'd161;
		data_a[3952]<=8'd170;
		data_a[3953]<=8'd174;
		data_a[3954]<=8'd158;
		data_a[3955]<=8'd178;
		data_a[3956]<=8'd207;
		data_a[3957]<=8'd228;
		data_a[3958]<=8'd223;
		data_a[3959]<=8'd226;
		data_a[3960]<=8'd226;
		data_a[3961]<=8'd228;
		data_a[3962]<=8'd216;
		data_a[3963]<=8'd231;
		data_a[3964]<=8'd223;
		data_a[3965]<=8'd224;
		data_a[3966]<=8'd222;
		data_a[3967]<=8'd219;
		data_a[3968]<=8'd221;
		data_a[3969]<=8'd225;
		data_a[3970]<=8'd210;
		data_a[3971]<=8'd212;
		data_a[3972]<=8'd218;
		data_a[3973]<=8'd217;
		data_a[3974]<=8'd216;
		data_a[3975]<=8'd216;
		data_a[3976]<=8'd217;
		data_a[3977]<=8'd213;
		data_a[3978]<=8'd158;
		data_a[3979]<=8'd121;
		data_a[3980]<=8'd119;
		data_a[3981]<=8'd116;
		data_a[3982]<=8'd126;
		data_a[3983]<=8'd137;
		data_a[3984]<=8'd97;
		data_a[3985]<=8'd98;
		data_a[3986]<=8'd104;
		data_a[3987]<=8'd93;
		data_a[3988]<=8'd104;
		data_a[3989]<=8'd91;
		data_a[3990]<=8'd82;
		data_a[3991]<=8'd75;
		data_a[3992]<=8'd76;
		data_a[3993]<=8'd68;
		data_a[3994]<=8'd69;
		data_a[3995]<=8'd70;
		data_a[3996]<=8'd76;
		data_a[3997]<=8'd76;
		data_a[3998]<=8'd73;
		data_a[3999]<=8'd71;
		data_a[4000]<=8'd79;
		data_a[4001]<=8'd82;
		data_a[4002]<=8'd90;
		data_a[4003]<=8'd92;
		data_a[4004]<=8'd94;
		data_a[4005]<=8'd96;
		data_a[4006]<=8'd95;
		data_a[4007]<=8'd92;
		data_a[4008]<=8'd92;
		data_a[4009]<=8'd91;
		data_a[4010]<=8'd91;
		data_a[4011]<=8'd93;
		data_a[4012]<=8'd96;
		data_a[4013]<=8'd97;
		data_a[4014]<=8'd94;
		data_a[4015]<=8'd95;
		data_a[4016]<=8'd96;
		data_a[4017]<=8'd103;
		data_a[4018]<=8'd104;
		data_a[4019]<=8'd116;
		data_a[4020]<=8'd115;
		data_a[4021]<=8'd139;
		data_a[4022]<=8'd163;
		data_a[4023]<=8'd162;
		data_a[4024]<=8'd201;
		data_a[4025]<=8'd211;
		data_a[4026]<=8'd218;
		data_a[4027]<=8'd220;
		data_a[4028]<=8'd216;
		data_a[4029]<=8'd223;
		data_a[4030]<=8'd224;
		data_a[4031]<=8'd231;
		data_a[4032]<=8'd233;
		data_a[4033]<=8'd234;
		data_a[4034]<=8'd253;
		data_a[4035]<=8'd254;
		data_a[4036]<=8'd249;
		data_a[4037]<=8'd245;
		data_a[4038]<=8'd239;
		data_a[4039]<=8'd243;
		data_a[4040]<=8'd243;
		data_a[4041]<=8'd247;
		data_a[4042]<=8'd241;
		data_a[4043]<=8'd238;
		data_a[4044]<=8'd238;
		data_a[4045]<=8'd238;
		data_a[4046]<=8'd236;
		data_a[4047]<=8'd234;
		data_a[4048]<=8'd231;
		data_a[4049]<=8'd230;
		data_a[4050]<=8'd254;
		data_a[4051]<=8'd187;
		data_a[4052]<=8'd175;
		data_a[4053]<=8'd176;
		data_a[4054]<=8'd140;
		data_a[4055]<=8'd114;
		data_a[4056]<=8'd128;
		data_a[4057]<=8'd148;
		data_a[4058]<=8'd204;
		data_a[4059]<=8'd209;
		data_a[4060]<=8'd214;
		data_a[4061]<=8'd211;
		data_a[4062]<=8'd220;
		data_a[4063]<=8'd214;
		data_a[4064]<=8'd209;
		data_a[4065]<=8'd212;
		data_a[4066]<=8'd215;
		data_a[4067]<=8'd210;
		data_a[4068]<=8'd211;
		data_a[4069]<=8'd216;
		data_a[4070]<=8'd216;
		data_a[4071]<=8'd193;
		data_a[4072]<=8'd217;
		data_a[4073]<=8'd212;
		data_a[4074]<=8'd217;
		data_a[4075]<=8'd213;
		data_a[4076]<=8'd212;
		data_a[4077]<=8'd210;
		data_a[4078]<=8'd210;
		data_a[4079]<=8'd212;
		data_a[4080]<=8'd213;
		data_a[4081]<=8'd210;
		data_a[4082]<=8'd208;
		data_a[4083]<=8'd179;
		data_a[4084]<=8'd182;
		data_a[4085]<=8'd138;
		data_a[4086]<=8'd168;
		data_a[4087]<=8'd154;
		data_a[4088]<=8'd127;
		data_a[4089]<=8'd120;
		data_a[4090]<=8'd127;
		data_a[4091]<=8'd124;
		data_a[4092]<=8'd111;
		data_a[4093]<=8'd112;
		data_a[4094]<=8'd100;
		data_a[4095]<=8'd122;
		data_a[4096]<=8'd98;
		data_a[4097]<=8'd110;
		data_a[4098]<=8'd172;
		data_a[4099]<=8'd156;
		data_a[4100]<=8'd151;
		data_a[4101]<=8'd182;
		data_a[4102]<=8'd157;
		data_a[4103]<=8'd176;
		data_a[4104]<=8'd171;
		data_a[4105]<=8'd156;
		data_a[4106]<=8'd202;
		data_a[4107]<=8'd195;
		data_a[4108]<=8'd182;
		data_a[4109]<=8'd170;
		data_a[4110]<=8'd207;
		data_a[4111]<=8'd223;
		data_a[4112]<=8'd225;
		data_a[4113]<=8'd215;
		data_a[4114]<=8'd225;
		data_a[4115]<=8'd226;
		data_a[4116]<=8'd222;
		data_a[4117]<=8'd214;
		data_a[4118]<=8'd210;
		data_a[4119]<=8'd215;
		data_a[4120]<=8'd212;
		data_a[4121]<=8'd219;
		data_a[4122]<=8'd222;
		data_a[4123]<=8'd211;
		data_a[4124]<=8'd219;
		data_a[4125]<=8'd218;
		data_a[4126]<=8'd213;
		data_a[4127]<=8'd215;
		data_a[4128]<=8'd116;
		data_a[4129]<=8'd108;
		data_a[4130]<=8'd117;
		data_a[4131]<=8'd101;
		data_a[4132]<=8'd126;
		data_a[4133]<=8'd75;
		data_a[4134]<=8'd86;
		data_a[4135]<=8'd106;
		data_a[4136]<=8'd74;
		data_a[4137]<=8'd117;
		data_a[4138]<=8'd89;
		data_a[4139]<=8'd87;
		data_a[4140]<=8'd82;
		data_a[4141]<=8'd72;
		data_a[4142]<=8'd71;
		data_a[4143]<=8'd71;
		data_a[4144]<=8'd74;
		data_a[4145]<=8'd73;
		data_a[4146]<=8'd73;
		data_a[4147]<=8'd78;
		data_a[4148]<=8'd81;
		data_a[4149]<=8'd84;
		data_a[4150]<=8'd94;
		data_a[4151]<=8'd95;
		data_a[4152]<=8'd101;
		data_a[4153]<=8'd100;
		data_a[4154]<=8'd103;
		data_a[4155]<=8'd107;
		data_a[4156]<=8'd108;
		data_a[4157]<=8'd107;
		data_a[4158]<=8'd107;
		data_a[4159]<=8'd104;
		data_a[4160]<=8'd100;
		data_a[4161]<=8'd100;
		data_a[4162]<=8'd96;
		data_a[4163]<=8'd98;
		data_a[4164]<=8'd97;
		data_a[4165]<=8'd98;
		data_a[4166]<=8'd99;
		data_a[4167]<=8'd102;
		data_a[4168]<=8'd101;
		data_a[4169]<=8'd105;
		data_a[4170]<=8'd117;
		data_a[4171]<=8'd126;
		data_a[4172]<=8'd135;
		data_a[4173]<=8'd132;
		data_a[4174]<=8'd222;
		data_a[4175]<=8'd218;
		data_a[4176]<=8'd220;
		data_a[4177]<=8'd218;
		data_a[4178]<=8'd223;
		data_a[4179]<=8'd224;
		data_a[4180]<=8'd225;
		data_a[4181]<=8'd227;
		data_a[4182]<=8'd230;
		data_a[4183]<=8'd224;
		data_a[4184]<=8'd233;
		data_a[4185]<=8'd229;
		data_a[4186]<=8'd241;
		data_a[4187]<=8'd240;
		data_a[4188]<=8'd238;
		data_a[4189]<=8'd240;
		data_a[4190]<=8'd239;
		data_a[4191]<=8'd241;
		data_a[4192]<=8'd239;
		data_a[4193]<=8'd238;
		data_a[4194]<=8'd236;
		data_a[4195]<=8'd235;
		data_a[4196]<=8'd234;
		data_a[4197]<=8'd232;
		data_a[4198]<=8'd230;
		data_a[4199]<=8'd230;
		data_a[4200]<=8'd254;
		data_a[4201]<=8'd213;
		data_a[4202]<=8'd187;
		data_a[4203]<=8'd159;
		data_a[4204]<=8'd167;
		data_a[4205]<=8'd151;
		data_a[4206]<=8'd114;
		data_a[4207]<=8'd126;
		data_a[4208]<=8'd178;
		data_a[4209]<=8'd212;
		data_a[4210]<=8'd205;
		data_a[4211]<=8'd216;
		data_a[4212]<=8'd207;
		data_a[4213]<=8'd211;
		data_a[4214]<=8'd215;
		data_a[4215]<=8'd213;
		data_a[4216]<=8'd215;
		data_a[4217]<=8'd210;
		data_a[4218]<=8'd213;
		data_a[4219]<=8'd212;
		data_a[4220]<=8'd210;
		data_a[4221]<=8'd216;
		data_a[4222]<=8'd195;
		data_a[4223]<=8'd211;
		data_a[4224]<=8'd211;
		data_a[4225]<=8'd207;
		data_a[4226]<=8'd207;
		data_a[4227]<=8'd215;
		data_a[4228]<=8'd214;
		data_a[4229]<=8'd210;
		data_a[4230]<=8'd205;
		data_a[4231]<=8'd206;
		data_a[4232]<=8'd191;
		data_a[4233]<=8'd179;
		data_a[4234]<=8'd175;
		data_a[4235]<=8'd125;
		data_a[4236]<=8'd134;
		data_a[4237]<=8'd138;
		data_a[4238]<=8'd116;
		data_a[4239]<=8'd104;
		data_a[4240]<=8'd132;
		data_a[4241]<=8'd122;
		data_a[4242]<=8'd98;
		data_a[4243]<=8'd97;
		data_a[4244]<=8'd105;
		data_a[4245]<=8'd106;
		data_a[4246]<=8'd103;
		data_a[4247]<=8'd108;
		data_a[4248]<=8'd131;
		data_a[4249]<=8'd145;
		data_a[4250]<=8'd144;
		data_a[4251]<=8'd145;
		data_a[4252]<=8'd141;
		data_a[4253]<=8'd144;
		data_a[4254]<=8'd197;
		data_a[4255]<=8'd153;
		data_a[4256]<=8'd146;
		data_a[4257]<=8'd178;
		data_a[4258]<=8'd170;
		data_a[4259]<=8'd162;
		data_a[4260]<=8'd153;
		data_a[4261]<=8'd185;
		data_a[4262]<=8'd225;
		data_a[4263]<=8'd225;
		data_a[4264]<=8'd220;
		data_a[4265]<=8'd223;
		data_a[4266]<=8'd225;
		data_a[4267]<=8'd222;
		data_a[4268]<=8'd217;
		data_a[4269]<=8'd213;
		data_a[4270]<=8'd219;
		data_a[4271]<=8'd215;
		data_a[4272]<=8'd215;
		data_a[4273]<=8'd218;
		data_a[4274]<=8'd212;
		data_a[4275]<=8'd219;
		data_a[4276]<=8'd214;
		data_a[4277]<=8'd222;
		data_a[4278]<=8'd105;
		data_a[4279]<=8'd129;
		data_a[4280]<=8'd110;
		data_a[4281]<=8'd108;
		data_a[4282]<=8'd90;
		data_a[4283]<=8'd84;
		data_a[4284]<=8'd89;
		data_a[4285]<=8'd98;
		data_a[4286]<=8'd110;
		data_a[4287]<=8'd98;
		data_a[4288]<=8'd89;
		data_a[4289]<=8'd82;
		data_a[4290]<=8'd70;
		data_a[4291]<=8'd67;
		data_a[4292]<=8'd68;
		data_a[4293]<=8'd74;
		data_a[4294]<=8'd71;
		data_a[4295]<=8'd67;
		data_a[4296]<=8'd74;
		data_a[4297]<=8'd82;
		data_a[4298]<=8'd89;
		data_a[4299]<=8'd95;
		data_a[4300]<=8'd106;
		data_a[4301]<=8'd107;
		data_a[4302]<=8'd111;
		data_a[4303]<=8'd111;
		data_a[4304]<=8'd114;
		data_a[4305]<=8'd117;
		data_a[4306]<=8'd116;
		data_a[4307]<=8'd115;
		data_a[4308]<=8'd116;
		data_a[4309]<=8'd117;
		data_a[4310]<=8'd116;
		data_a[4311]<=8'd117;
		data_a[4312]<=8'd110;
		data_a[4313]<=8'd105;
		data_a[4314]<=8'd102;
		data_a[4315]<=8'd95;
		data_a[4316]<=8'd94;
		data_a[4317]<=8'd95;
		data_a[4318]<=8'd101;
		data_a[4319]<=8'd99;
		data_a[4320]<=8'd121;
		data_a[4321]<=8'd136;
		data_a[4322]<=8'd136;
		data_a[4323]<=8'd141;
		data_a[4324]<=8'd214;
		data_a[4325]<=8'd221;
		data_a[4326]<=8'd217;
		data_a[4327]<=8'd221;
		data_a[4328]<=8'd221;
		data_a[4329]<=8'd217;
		data_a[4330]<=8'd222;
		data_a[4331]<=8'd223;
		data_a[4332]<=8'd229;
		data_a[4333]<=8'd230;
		data_a[4334]<=8'd234;
		data_a[4335]<=8'd233;
		data_a[4336]<=8'd237;
		data_a[4337]<=8'd237;
		data_a[4338]<=8'd240;
		data_a[4339]<=8'd238;
		data_a[4340]<=8'd239;
		data_a[4341]<=8'd236;
		data_a[4342]<=8'd237;
		data_a[4343]<=8'd236;
		data_a[4344]<=8'd234;
		data_a[4345]<=8'd233;
		data_a[4346]<=8'd232;
		data_a[4347]<=8'd231;
		data_a[4348]<=8'd230;
		data_a[4349]<=8'd230;
		data_a[4350]<=8'd254;
		data_a[4351]<=8'd208;
		data_a[4352]<=8'd179;
		data_a[4353]<=8'd181;
		data_a[4354]<=8'd172;
		data_a[4355]<=8'd186;
		data_a[4356]<=8'd163;
		data_a[4357]<=8'd124;
		data_a[4358]<=8'd187;
		data_a[4359]<=8'd157;
		data_a[4360]<=8'd156;
		data_a[4361]<=8'd204;
		data_a[4362]<=8'd215;
		data_a[4363]<=8'd217;
		data_a[4364]<=8'd219;
		data_a[4365]<=8'd207;
		data_a[4366]<=8'd211;
		data_a[4367]<=8'd212;
		data_a[4368]<=8'd214;
		data_a[4369]<=8'd213;
		data_a[4370]<=8'd189;
		data_a[4371]<=8'd195;
		data_a[4372]<=8'd210;
		data_a[4373]<=8'd203;
		data_a[4374]<=8'd214;
		data_a[4375]<=8'd215;
		data_a[4376]<=8'd207;
		data_a[4377]<=8'd210;
		data_a[4378]<=8'd209;
		data_a[4379]<=8'd213;
		data_a[4380]<=8'd206;
		data_a[4381]<=8'd207;
		data_a[4382]<=8'd189;
		data_a[4383]<=8'd174;
		data_a[4384]<=8'd180;
		data_a[4385]<=8'd107;
		data_a[4386]<=8'd135;
		data_a[4387]<=8'd173;
		data_a[4388]<=8'd106;
		data_a[4389]<=8'd104;
		data_a[4390]<=8'd110;
		data_a[4391]<=8'd107;
		data_a[4392]<=8'd89;
		data_a[4393]<=8'd90;
		data_a[4394]<=8'd108;
		data_a[4395]<=8'd112;
		data_a[4396]<=8'd97;
		data_a[4397]<=8'd110;
		data_a[4398]<=8'd139;
		data_a[4399]<=8'd127;
		data_a[4400]<=8'd123;
		data_a[4401]<=8'd138;
		data_a[4402]<=8'd128;
		data_a[4403]<=8'd124;
		data_a[4404]<=8'd140;
		data_a[4405]<=8'd131;
		data_a[4406]<=8'd137;
		data_a[4407]<=8'd168;
		data_a[4408]<=8'd168;
		data_a[4409]<=8'd151;
		data_a[4410]<=8'd172;
		data_a[4411]<=8'd136;
		data_a[4412]<=8'd218;
		data_a[4413]<=8'd228;
		data_a[4414]<=8'd225;
		data_a[4415]<=8'd222;
		data_a[4416]<=8'd219;
		data_a[4417]<=8'd219;
		data_a[4418]<=8'd217;
		data_a[4419]<=8'd213;
		data_a[4420]<=8'd224;
		data_a[4421]<=8'd217;
		data_a[4422]<=8'd216;
		data_a[4423]<=8'd220;
		data_a[4424]<=8'd218;
		data_a[4425]<=8'd214;
		data_a[4426]<=8'd224;
		data_a[4427]<=8'd203;
		data_a[4428]<=8'd145;
		data_a[4429]<=8'd114;
		data_a[4430]<=8'd106;
		data_a[4431]<=8'd97;
		data_a[4432]<=8'd90;
		data_a[4433]<=8'd106;
		data_a[4434]<=8'd106;
		data_a[4435]<=8'd97;
		data_a[4436]<=8'd101;
		data_a[4437]<=8'd86;
		data_a[4438]<=8'd87;
		data_a[4439]<=8'd76;
		data_a[4440]<=8'd67;
		data_a[4441]<=8'd73;
		data_a[4442]<=8'd71;
		data_a[4443]<=8'd73;
		data_a[4444]<=8'd74;
		data_a[4445]<=8'd83;
		data_a[4446]<=8'd84;
		data_a[4447]<=8'd92;
		data_a[4448]<=8'd100;
		data_a[4449]<=8'd105;
		data_a[4450]<=8'd115;
		data_a[4451]<=8'd116;
		data_a[4452]<=8'd124;
		data_a[4453]<=8'd125;
		data_a[4454]<=8'd127;
		data_a[4455]<=8'd130;
		data_a[4456]<=8'd128;
		data_a[4457]<=8'd126;
		data_a[4458]<=8'd129;
		data_a[4459]<=8'd132;
		data_a[4460]<=8'd132;
		data_a[4461]<=8'd133;
		data_a[4462]<=8'd128;
		data_a[4463]<=8'd122;
		data_a[4464]<=8'd114;
		data_a[4465]<=8'd101;
		data_a[4466]<=8'd95;
		data_a[4467]<=8'd95;
		data_a[4468]<=8'd105;
		data_a[4469]<=8'd102;
		data_a[4470]<=8'd103;
		data_a[4471]<=8'd117;
		data_a[4472]<=8'd125;
		data_a[4473]<=8'd142;
		data_a[4474]<=8'd223;
		data_a[4475]<=8'd217;
		data_a[4476]<=8'd214;
		data_a[4477]<=8'd220;
		data_a[4478]<=8'd224;
		data_a[4479]<=8'd220;
		data_a[4480]<=8'd227;
		data_a[4481]<=8'd228;
		data_a[4482]<=8'd231;
		data_a[4483]<=8'd233;
		data_a[4484]<=8'd233;
		data_a[4485]<=8'd235;
		data_a[4486]<=8'd235;
		data_a[4487]<=8'd233;
		data_a[4488]<=8'd235;
		data_a[4489]<=8'd234;
		data_a[4490]<=8'd240;
		data_a[4491]<=8'd237;
		data_a[4492]<=8'd237;
		data_a[4493]<=8'd233;
		data_a[4494]<=8'd233;
		data_a[4495]<=8'd232;
		data_a[4496]<=8'd230;
		data_a[4497]<=8'd230;
		data_a[4498]<=8'd230;
		data_a[4499]<=8'd230;
		data_a[4500]<=8'd252;
		data_a[4501]<=8'd199;
		data_a[4502]<=8'd173;
		data_a[4503]<=8'd171;
		data_a[4504]<=8'd163;
		data_a[4505]<=8'd142;
		data_a[4506]<=8'd183;
		data_a[4507]<=8'd129;
		data_a[4508]<=8'd201;
		data_a[4509]<=8'd135;
		data_a[4510]<=8'd128;
		data_a[4511]<=8'd211;
		data_a[4512]<=8'd209;
		data_a[4513]<=8'd211;
		data_a[4514]<=8'd221;
		data_a[4515]<=8'd214;
		data_a[4516]<=8'd215;
		data_a[4517]<=8'd209;
		data_a[4518]<=8'd190;
		data_a[4519]<=8'd195;
		data_a[4520]<=8'd218;
		data_a[4521]<=8'd213;
		data_a[4522]<=8'd206;
		data_a[4523]<=8'd210;
		data_a[4524]<=8'd200;
		data_a[4525]<=8'd205;
		data_a[4526]<=8'd208;
		data_a[4527]<=8'd207;
		data_a[4528]<=8'd214;
		data_a[4529]<=8'd196;
		data_a[4530]<=8'd175;
		data_a[4531]<=8'd163;
		data_a[4532]<=8'd168;
		data_a[4533]<=8'd181;
		data_a[4534]<=8'd153;
		data_a[4535]<=8'd113;
		data_a[4536]<=8'd92;
		data_a[4537]<=8'd102;
		data_a[4538]<=8'd97;
		data_a[4539]<=8'd90;
		data_a[4540]<=8'd92;
		data_a[4541]<=8'd91;
		data_a[4542]<=8'd87;
		data_a[4543]<=8'd83;
		data_a[4544]<=8'd104;
		data_a[4545]<=8'd90;
		data_a[4546]<=8'd95;
		data_a[4547]<=8'd108;
		data_a[4548]<=8'd110;
		data_a[4549]<=8'd121;
		data_a[4550]<=8'd120;
		data_a[4551]<=8'd137;
		data_a[4552]<=8'd132;
		data_a[4553]<=8'd125;
		data_a[4554]<=8'd135;
		data_a[4555]<=8'd128;
		data_a[4556]<=8'd125;
		data_a[4557]<=8'd149;
		data_a[4558]<=8'd193;
		data_a[4559]<=8'd197;
		data_a[4560]<=8'd157;
		data_a[4561]<=8'd159;
		data_a[4562]<=8'd143;
		data_a[4563]<=8'd221;
		data_a[4564]<=8'd217;
		data_a[4565]<=8'd219;
		data_a[4566]<=8'd223;
		data_a[4567]<=8'd223;
		data_a[4568]<=8'd218;
		data_a[4569]<=8'd212;
		data_a[4570]<=8'd215;
		data_a[4571]<=8'd218;
		data_a[4572]<=8'd214;
		data_a[4573]<=8'd215;
		data_a[4574]<=8'd221;
		data_a[4575]<=8'd212;
		data_a[4576]<=8'd210;
		data_a[4577]<=8'd208;
		data_a[4578]<=8'd118;
		data_a[4579]<=8'd109;
		data_a[4580]<=8'd112;
		data_a[4581]<=8'd109;
		data_a[4582]<=8'd94;
		data_a[4583]<=8'd115;
		data_a[4584]<=8'd100;
		data_a[4585]<=8'd102;
		data_a[4586]<=8'd90;
		data_a[4587]<=8'd91;
		data_a[4588]<=8'd67;
		data_a[4589]<=8'd68;
		data_a[4590]<=8'd69;
		data_a[4591]<=8'd74;
		data_a[4592]<=8'd78;
		data_a[4593]<=8'd84;
		data_a[4594]<=8'd86;
		data_a[4595]<=8'd87;
		data_a[4596]<=8'd95;
		data_a[4597]<=8'd107;
		data_a[4598]<=8'd118;
		data_a[4599]<=8'd125;
		data_a[4600]<=8'd133;
		data_a[4601]<=8'd131;
		data_a[4602]<=8'd135;
		data_a[4603]<=8'd134;
		data_a[4604]<=8'd139;
		data_a[4605]<=8'd142;
		data_a[4606]<=8'd142;
		data_a[4607]<=8'd143;
		data_a[4608]<=8'd147;
		data_a[4609]<=8'd149;
		data_a[4610]<=8'd147;
		data_a[4611]<=8'd146;
		data_a[4612]<=8'd147;
		data_a[4613]<=8'd149;
		data_a[4614]<=8'd137;
		data_a[4615]<=8'd120;
		data_a[4616]<=8'd109;
		data_a[4617]<=8'd103;
		data_a[4618]<=8'd107;
		data_a[4619]<=8'd107;
		data_a[4620]<=8'd111;
		data_a[4621]<=8'd110;
		data_a[4622]<=8'd116;
		data_a[4623]<=8'd172;
		data_a[4624]<=8'd213;
		data_a[4625]<=8'd214;
		data_a[4626]<=8'd220;
		data_a[4627]<=8'd217;
		data_a[4628]<=8'd219;
		data_a[4629]<=8'd219;
		data_a[4630]<=8'd222;
		data_a[4631]<=8'd230;
		data_a[4632]<=8'd229;
		data_a[4633]<=8'd229;
		data_a[4634]<=8'd230;
		data_a[4635]<=8'd229;
		data_a[4636]<=8'd232;
		data_a[4637]<=8'd236;
		data_a[4638]<=8'd239;
		data_a[4639]<=8'd237;
		data_a[4640]<=8'd233;
		data_a[4641]<=8'd229;
		data_a[4642]<=8'd231;
		data_a[4643]<=8'd233;
		data_a[4644]<=8'd232;
		data_a[4645]<=8'd232;
		data_a[4646]<=8'd230;
		data_a[4647]<=8'd229;
		data_a[4648]<=8'd229;
		data_a[4649]<=8'd228;
		data_a[4650]<=8'd254;
		data_a[4651]<=8'd185;
		data_a[4652]<=8'd167;
		data_a[4653]<=8'd164;
		data_a[4654]<=8'd167;
		data_a[4655]<=8'd185;
		data_a[4656]<=8'd124;
		data_a[4657]<=8'd141;
		data_a[4658]<=8'd201;
		data_a[4659]<=8'd108;
		data_a[4660]<=8'd188;
		data_a[4661]<=8'd123;
		data_a[4662]<=8'd153;
		data_a[4663]<=8'd202;
		data_a[4664]<=8'd207;
		data_a[4665]<=8'd198;
		data_a[4666]<=8'd191;
		data_a[4667]<=8'd202;
		data_a[4668]<=8'd217;
		data_a[4669]<=8'd212;
		data_a[4670]<=8'd209;
		data_a[4671]<=8'd211;
		data_a[4672]<=8'd210;
		data_a[4673]<=8'd208;
		data_a[4674]<=8'd210;
		data_a[4675]<=8'd195;
		data_a[4676]<=8'd202;
		data_a[4677]<=8'd195;
		data_a[4678]<=8'd213;
		data_a[4679]<=8'd161;
		data_a[4680]<=8'd141;
		data_a[4681]<=8'd132;
		data_a[4682]<=8'd127;
		data_a[4683]<=8'd124;
		data_a[4684]<=8'd142;
		data_a[4685]<=8'd120;
		data_a[4686]<=8'd102;
		data_a[4687]<=8'd92;
		data_a[4688]<=8'd82;
		data_a[4689]<=8'd89;
		data_a[4690]<=8'd81;
		data_a[4691]<=8'd84;
		data_a[4692]<=8'd78;
		data_a[4693]<=8'd85;
		data_a[4694]<=8'd86;
		data_a[4695]<=8'd82;
		data_a[4696]<=8'd92;
		data_a[4697]<=8'd92;
		data_a[4698]<=8'd86;
		data_a[4699]<=8'd117;
		data_a[4700]<=8'd118;
		data_a[4701]<=8'd124;
		data_a[4702]<=8'd122;
		data_a[4703]<=8'd119;
		data_a[4704]<=8'd117;
		data_a[4705]<=8'd117;
		data_a[4706]<=8'd117;
		data_a[4707]<=8'd127;
		data_a[4708]<=8'd180;
		data_a[4709]<=8'd176;
		data_a[4710]<=8'd118;
		data_a[4711]<=8'd152;
		data_a[4712]<=8'd123;
		data_a[4713]<=8'd168;
		data_a[4714]<=8'd222;
		data_a[4715]<=8'd220;
		data_a[4716]<=8'd217;
		data_a[4717]<=8'd217;
		data_a[4718]<=8'd217;
		data_a[4719]<=8'd218;
		data_a[4720]<=8'd210;
		data_a[4721]<=8'd219;
		data_a[4722]<=8'd216;
		data_a[4723]<=8'd217;
		data_a[4724]<=8'd211;
		data_a[4725]<=8'd216;
		data_a[4726]<=8'd212;
		data_a[4727]<=8'd160;
		data_a[4728]<=8'd103;
		data_a[4729]<=8'd103;
		data_a[4730]<=8'd105;
		data_a[4731]<=8'd111;
		data_a[4732]<=8'd132;
		data_a[4733]<=8'd116;
		data_a[4734]<=8'd96;
		data_a[4735]<=8'd87;
		data_a[4736]<=8'd91;
		data_a[4737]<=8'd62;
		data_a[4738]<=8'd73;
		data_a[4739]<=8'd68;
		data_a[4740]<=8'd75;
		data_a[4741]<=8'd83;
		data_a[4742]<=8'd91;
		data_a[4743]<=8'd88;
		data_a[4744]<=8'd97;
		data_a[4745]<=8'd108;
		data_a[4746]<=8'd110;
		data_a[4747]<=8'd121;
		data_a[4748]<=8'd131;
		data_a[4749]<=8'd136;
		data_a[4750]<=8'd143;
		data_a[4751]<=8'd140;
		data_a[4752]<=8'd146;
		data_a[4753]<=8'd147;
		data_a[4754]<=8'd146;
		data_a[4755]<=8'd149;
		data_a[4756]<=8'd150;
		data_a[4757]<=8'd152;
		data_a[4758]<=8'd158;
		data_a[4759]<=8'd162;
		data_a[4760]<=8'd160;
		data_a[4761]<=8'd158;
		data_a[4762]<=8'd163;
		data_a[4763]<=8'd174;
		data_a[4764]<=8'd155;
		data_a[4765]<=8'd135;
		data_a[4766]<=8'd119;
		data_a[4767]<=8'd108;
		data_a[4768]<=8'd104;
		data_a[4769]<=8'd109;
		data_a[4770]<=8'd105;
		data_a[4771]<=8'd119;
		data_a[4772]<=8'd116;
		data_a[4773]<=8'd175;
		data_a[4774]<=8'd220;
		data_a[4775]<=8'd217;
		data_a[4776]<=8'd222;
		data_a[4777]<=8'd216;
		data_a[4778]<=8'd220;
		data_a[4779]<=8'd222;
		data_a[4780]<=8'd217;
		data_a[4781]<=8'd230;
		data_a[4782]<=8'd229;
		data_a[4783]<=8'd228;
		data_a[4784]<=8'd233;
		data_a[4785]<=8'd229;
		data_a[4786]<=8'd232;
		data_a[4787]<=8'd233;
		data_a[4788]<=8'd231;
		data_a[4789]<=8'd235;
		data_a[4790]<=8'd232;
		data_a[4791]<=8'd234;
		data_a[4792]<=8'd232;
		data_a[4793]<=8'd232;
		data_a[4794]<=8'd232;
		data_a[4795]<=8'd232;
		data_a[4796]<=8'd231;
		data_a[4797]<=8'd230;
		data_a[4798]<=8'd228;
		data_a[4799]<=8'd227;
		data_a[4800]<=8'd253;
		data_a[4801]<=8'd204;
		data_a[4802]<=8'd222;
		data_a[4803]<=8'd189;
		data_a[4804]<=8'd198;
		data_a[4805]<=8'd179;
		data_a[4806]<=8'd131;
		data_a[4807]<=8'd113;
		data_a[4808]<=8'd182;
		data_a[4809]<=8'd131;
		data_a[4810]<=8'd186;
		data_a[4811]<=8'd171;
		data_a[4812]<=8'd206;
		data_a[4813]<=8'd201;
		data_a[4814]<=8'd192;
		data_a[4815]<=8'd208;
		data_a[4816]<=8'd210;
		data_a[4817]<=8'd210;
		data_a[4818]<=8'd207;
		data_a[4819]<=8'd213;
		data_a[4820]<=8'd210;
		data_a[4821]<=8'd208;
		data_a[4822]<=8'd215;
		data_a[4823]<=8'd205;
		data_a[4824]<=8'd213;
		data_a[4825]<=8'd208;
		data_a[4826]<=8'd198;
		data_a[4827]<=8'd188;
		data_a[4828]<=8'd108;
		data_a[4829]<=8'd134;
		data_a[4830]<=8'd141;
		data_a[4831]<=8'd115;
		data_a[4832]<=8'd121;
		data_a[4833]<=8'd119;
		data_a[4834]<=8'd104;
		data_a[4835]<=8'd118;
		data_a[4836]<=8'd111;
		data_a[4837]<=8'd85;
		data_a[4838]<=8'd83;
		data_a[4839]<=8'd84;
		data_a[4840]<=8'd81;
		data_a[4841]<=8'd85;
		data_a[4842]<=8'd83;
		data_a[4843]<=8'd88;
		data_a[4844]<=8'd79;
		data_a[4845]<=8'd79;
		data_a[4846]<=8'd87;
		data_a[4847]<=8'd92;
		data_a[4848]<=8'd93;
		data_a[4849]<=8'd107;
		data_a[4850]<=8'd110;
		data_a[4851]<=8'd122;
		data_a[4852]<=8'd119;
		data_a[4853]<=8'd118;
		data_a[4854]<=8'd120;
		data_a[4855]<=8'd110;
		data_a[4856]<=8'd115;
		data_a[4857]<=8'd111;
		data_a[4858]<=8'd166;
		data_a[4859]<=8'd166;
		data_a[4860]<=8'd135;
		data_a[4861]<=8'd149;
		data_a[4862]<=8'd117;
		data_a[4863]<=8'd131;
		data_a[4864]<=8'd228;
		data_a[4865]<=8'd218;
		data_a[4866]<=8'd219;
		data_a[4867]<=8'd218;
		data_a[4868]<=8'd217;
		data_a[4869]<=8'd218;
		data_a[4870]<=8'd217;
		data_a[4871]<=8'd212;
		data_a[4872]<=8'd216;
		data_a[4873]<=8'd216;
		data_a[4874]<=8'd215;
		data_a[4875]<=8'd213;
		data_a[4876]<=8'd218;
		data_a[4877]<=8'd100;
		data_a[4878]<=8'd111;
		data_a[4879]<=8'd105;
		data_a[4880]<=8'd127;
		data_a[4881]<=8'd116;
		data_a[4882]<=8'd107;
		data_a[4883]<=8'd102;
		data_a[4884]<=8'd97;
		data_a[4885]<=8'd85;
		data_a[4886]<=8'd63;
		data_a[4887]<=8'd73;
		data_a[4888]<=8'd67;
		data_a[4889]<=8'd69;
		data_a[4890]<=8'd79;
		data_a[4891]<=8'd88;
		data_a[4892]<=8'd95;
		data_a[4893]<=8'd97;
		data_a[4894]<=8'd101;
		data_a[4895]<=8'd113;
		data_a[4896]<=8'd126;
		data_a[4897]<=8'd134;
		data_a[4898]<=8'd142;
		data_a[4899]<=8'd148;
		data_a[4900]<=8'd154;
		data_a[4901]<=8'd154;
		data_a[4902]<=8'd150;
		data_a[4903]<=8'd147;
		data_a[4904]<=8'd150;
		data_a[4905]<=8'd154;
		data_a[4906]<=8'd158;
		data_a[4907]<=8'd163;
		data_a[4908]<=8'd167;
		data_a[4909]<=8'd171;
		data_a[4910]<=8'd170;
		data_a[4911]<=8'd167;
		data_a[4912]<=8'd174;
		data_a[4913]<=8'd174;
		data_a[4914]<=8'd164;
		data_a[4915]<=8'd147;
		data_a[4916]<=8'd129;
		data_a[4917]<=8'd122;
		data_a[4918]<=8'd98;
		data_a[4919]<=8'd108;
		data_a[4920]<=8'd111;
		data_a[4921]<=8'd118;
		data_a[4922]<=8'd138;
		data_a[4923]<=8'd159;
		data_a[4924]<=8'd212;
		data_a[4925]<=8'd216;
		data_a[4926]<=8'd216;
		data_a[4927]<=8'd217;
		data_a[4928]<=8'd219;
		data_a[4929]<=8'd221;
		data_a[4930]<=8'd220;
		data_a[4931]<=8'd224;
		data_a[4932]<=8'd224;
		data_a[4933]<=8'd231;
		data_a[4934]<=8'd229;
		data_a[4935]<=8'd229;
		data_a[4936]<=8'd232;
		data_a[4937]<=8'd230;
		data_a[4938]<=8'd231;
		data_a[4939]<=8'd233;
		data_a[4940]<=8'd234;
		data_a[4941]<=8'd231;
		data_a[4942]<=8'd230;
		data_a[4943]<=8'd231;
		data_a[4944]<=8'd230;
		data_a[4945]<=8'd231;
		data_a[4946]<=8'd231;
		data_a[4947]<=8'd230;
		data_a[4948]<=8'd228;
		data_a[4949]<=8'd225;
		data_a[4950]<=8'd254;
		data_a[4951]<=8'd197;
		data_a[4952]<=8'd197;
		data_a[4953]<=8'd136;
		data_a[4954]<=8'd124;
		data_a[4955]<=8'd160;
		data_a[4956]<=8'd212;
		data_a[4957]<=8'd140;
		data_a[4958]<=8'd114;
		data_a[4959]<=8'd216;
		data_a[4960]<=8'd195;
		data_a[4961]<=8'd196;
		data_a[4962]<=8'd201;
		data_a[4963]<=8'd204;
		data_a[4964]<=8'd222;
		data_a[4965]<=8'd206;
		data_a[4966]<=8'd210;
		data_a[4967]<=8'd210;
		data_a[4968]<=8'd208;
		data_a[4969]<=8'd211;
		data_a[4970]<=8'd210;
		data_a[4971]<=8'd209;
		data_a[4972]<=8'd213;
		data_a[4973]<=8'd207;
		data_a[4974]<=8'd209;
		data_a[4975]<=8'd203;
		data_a[4976]<=8'd199;
		data_a[4977]<=8'd111;
		data_a[4978]<=8'd178;
		data_a[4979]<=8'd200;
		data_a[4980]<=8'd128;
		data_a[4981]<=8'd102;
		data_a[4982]<=8'd109;
		data_a[4983]<=8'd117;
		data_a[4984]<=8'd111;
		data_a[4985]<=8'd107;
		data_a[4986]<=8'd93;
		data_a[4987]<=8'd93;
		data_a[4988]<=8'd80;
		data_a[4989]<=8'd80;
		data_a[4990]<=8'd83;
		data_a[4991]<=8'd80;
		data_a[4992]<=8'd75;
		data_a[4993]<=8'd79;
		data_a[4994]<=8'd77;
		data_a[4995]<=8'd82;
		data_a[4996]<=8'd84;
		data_a[4997]<=8'd85;
		data_a[4998]<=8'd87;
		data_a[4999]<=8'd100;
		data_a[5000]<=8'd107;
		data_a[5001]<=8'd115;
		data_a[5002]<=8'd114;
		data_a[5003]<=8'd123;
		data_a[5004]<=8'd113;
		data_a[5005]<=8'd113;
		data_a[5006]<=8'd112;
		data_a[5007]<=8'd110;
		data_a[5008]<=8'd152;
		data_a[5009]<=8'd164;
		data_a[5010]<=8'd143;
		data_a[5011]<=8'd139;
		data_a[5012]<=8'd109;
		data_a[5013]<=8'd126;
		data_a[5014]<=8'd184;
		data_a[5015]<=8'd220;
		data_a[5016]<=8'd214;
		data_a[5017]<=8'd215;
		data_a[5018]<=8'd220;
		data_a[5019]<=8'd214;
		data_a[5020]<=8'd222;
		data_a[5021]<=8'd215;
		data_a[5022]<=8'd211;
		data_a[5023]<=8'd216;
		data_a[5024]<=8'd214;
		data_a[5025]<=8'd218;
		data_a[5026]<=8'd202;
		data_a[5027]<=8'd108;
		data_a[5028]<=8'd97;
		data_a[5029]<=8'd104;
		data_a[5030]<=8'd114;
		data_a[5031]<=8'd97;
		data_a[5032]<=8'd101;
		data_a[5033]<=8'd96;
		data_a[5034]<=8'd86;
		data_a[5035]<=8'd69;
		data_a[5036]<=8'd70;
		data_a[5037]<=8'd66;
		data_a[5038]<=8'd72;
		data_a[5039]<=8'd75;
		data_a[5040]<=8'd85;
		data_a[5041]<=8'd94;
		data_a[5042]<=8'd102;
		data_a[5043]<=8'd107;
		data_a[5044]<=8'd114;
		data_a[5045]<=8'd127;
		data_a[5046]<=8'd138;
		data_a[5047]<=8'd149;
		data_a[5048]<=8'd157;
		data_a[5049]<=8'd160;
		data_a[5050]<=8'd161;
		data_a[5051]<=8'd160;
		data_a[5052]<=8'd159;
		data_a[5053]<=8'd161;
		data_a[5054]<=8'd160;
		data_a[5055]<=8'd162;
		data_a[5056]<=8'd168;
		data_a[5057]<=8'd173;
		data_a[5058]<=8'd177;
		data_a[5059]<=8'd176;
		data_a[5060]<=8'd174;
		data_a[5061]<=8'd173;
		data_a[5062]<=8'd179;
		data_a[5063]<=8'd171;
		data_a[5064]<=8'd169;
		data_a[5065]<=8'd168;
		data_a[5066]<=8'd149;
		data_a[5067]<=8'd135;
		data_a[5068]<=8'd113;
		data_a[5069]<=8'd101;
		data_a[5070]<=8'd109;
		data_a[5071]<=8'd121;
		data_a[5072]<=8'd140;
		data_a[5073]<=8'd146;
		data_a[5074]<=8'd218;
		data_a[5075]<=8'd217;
		data_a[5076]<=8'd218;
		data_a[5077]<=8'd217;
		data_a[5078]<=8'd219;
		data_a[5079]<=8'd220;
		data_a[5080]<=8'd220;
		data_a[5081]<=8'd223;
		data_a[5082]<=8'd225;
		data_a[5083]<=8'd229;
		data_a[5084]<=8'd229;
		data_a[5085]<=8'd229;
		data_a[5086]<=8'd232;
		data_a[5087]<=8'd231;
		data_a[5088]<=8'd231;
		data_a[5089]<=8'd233;
		data_a[5090]<=8'd233;
		data_a[5091]<=8'd232;
		data_a[5092]<=8'd231;
		data_a[5093]<=8'd233;
		data_a[5094]<=8'd232;
		data_a[5095]<=8'd232;
		data_a[5096]<=8'd232;
		data_a[5097]<=8'd230;
		data_a[5098]<=8'd228;
		data_a[5099]<=8'd226;
		data_a[5100]<=8'd254;
		data_a[5101]<=8'd208;
		data_a[5102]<=8'd202;
		data_a[5103]<=8'd151;
		data_a[5104]<=8'd212;
		data_a[5105]<=8'd211;
		data_a[5106]<=8'd116;
		data_a[5107]<=8'd179;
		data_a[5108]<=8'd194;
		data_a[5109]<=8'd192;
		data_a[5110]<=8'd201;
		data_a[5111]<=8'd205;
		data_a[5112]<=8'd215;
		data_a[5113]<=8'd205;
		data_a[5114]<=8'd220;
		data_a[5115]<=8'd208;
		data_a[5116]<=8'd211;
		data_a[5117]<=8'd211;
		data_a[5118]<=8'd210;
		data_a[5119]<=8'd210;
		data_a[5120]<=8'd210;
		data_a[5121]<=8'd210;
		data_a[5122]<=8'd209;
		data_a[5123]<=8'd206;
		data_a[5124]<=8'd206;
		data_a[5125]<=8'd211;
		data_a[5126]<=8'd187;
		data_a[5127]<=8'd172;
		data_a[5128]<=8'd165;
		data_a[5129]<=8'd179;
		data_a[5130]<=8'd120;
		data_a[5131]<=8'd110;
		data_a[5132]<=8'd109;
		data_a[5133]<=8'd141;
		data_a[5134]<=8'd117;
		data_a[5135]<=8'd107;
		data_a[5136]<=8'd88;
		data_a[5137]<=8'd91;
		data_a[5138]<=8'd83;
		data_a[5139]<=8'd77;
		data_a[5140]<=8'd74;
		data_a[5141]<=8'd74;
		data_a[5142]<=8'd76;
		data_a[5143]<=8'd79;
		data_a[5144]<=8'd76;
		data_a[5145]<=8'd81;
		data_a[5146]<=8'd80;
		data_a[5147]<=8'd81;
		data_a[5148]<=8'd94;
		data_a[5149]<=8'd105;
		data_a[5150]<=8'd106;
		data_a[5151]<=8'd117;
		data_a[5152]<=8'd121;
		data_a[5153]<=8'd131;
		data_a[5154]<=8'd114;
		data_a[5155]<=8'd112;
		data_a[5156]<=8'd107;
		data_a[5157]<=8'd98;
		data_a[5158]<=8'd133;
		data_a[5159]<=8'd138;
		data_a[5160]<=8'd134;
		data_a[5161]<=8'd132;
		data_a[5162]<=8'd115;
		data_a[5163]<=8'd110;
		data_a[5164]<=8'd127;
		data_a[5165]<=8'd214;
		data_a[5166]<=8'd218;
		data_a[5167]<=8'd215;
		data_a[5168]<=8'd216;
		data_a[5169]<=8'd214;
		data_a[5170]<=8'd207;
		data_a[5171]<=8'd198;
		data_a[5172]<=8'd207;
		data_a[5173]<=8'd216;
		data_a[5174]<=8'd213;
		data_a[5175]<=8'd210;
		data_a[5176]<=8'd218;
		data_a[5177]<=8'd114;
		data_a[5178]<=8'd95;
		data_a[5179]<=8'd112;
		data_a[5180]<=8'd110;
		data_a[5181]<=8'd99;
		data_a[5182]<=8'd83;
		data_a[5183]<=8'd99;
		data_a[5184]<=8'd66;
		data_a[5185]<=8'd75;
		data_a[5186]<=8'd75;
		data_a[5187]<=8'd79;
		data_a[5188]<=8'd78;
		data_a[5189]<=8'd83;
		data_a[5190]<=8'd93;
		data_a[5191]<=8'd102;
		data_a[5192]<=8'd111;
		data_a[5193]<=8'd119;
		data_a[5194]<=8'd128;
		data_a[5195]<=8'd141;
		data_a[5196]<=8'd151;
		data_a[5197]<=8'd161;
		data_a[5198]<=8'd168;
		data_a[5199]<=8'd168;
		data_a[5200]<=8'd167;
		data_a[5201]<=8'd166;
		data_a[5202]<=8'd167;
		data_a[5203]<=8'd170;
		data_a[5204]<=8'd172;
		data_a[5205]<=8'd172;
		data_a[5206]<=8'd176;
		data_a[5207]<=8'd180;
		data_a[5208]<=8'd181;
		data_a[5209]<=8'd179;
		data_a[5210]<=8'd178;
		data_a[5211]<=8'd180;
		data_a[5212]<=8'd187;
		data_a[5213]<=8'd178;
		data_a[5214]<=8'd173;
		data_a[5215]<=8'd173;
		data_a[5216]<=8'd160;
		data_a[5217]<=8'd147;
		data_a[5218]<=8'd134;
		data_a[5219]<=8'd112;
		data_a[5220]<=8'd109;
		data_a[5221]<=8'd112;
		data_a[5222]<=8'd138;
		data_a[5223]<=8'd164;
		data_a[5224]<=8'd214;
		data_a[5225]<=8'd215;
		data_a[5226]<=8'd216;
		data_a[5227]<=8'd223;
		data_a[5228]<=8'd219;
		data_a[5229]<=8'd219;
		data_a[5230]<=8'd221;
		data_a[5231]<=8'd222;
		data_a[5232]<=8'd226;
		data_a[5233]<=8'd227;
		data_a[5234]<=8'd229;
		data_a[5235]<=8'd228;
		data_a[5236]<=8'd230;
		data_a[5237]<=8'd229;
		data_a[5238]<=8'd229;
		data_a[5239]<=8'd230;
		data_a[5240]<=8'd231;
		data_a[5241]<=8'd231;
		data_a[5242]<=8'd231;
		data_a[5243]<=8'd232;
		data_a[5244]<=8'd232;
		data_a[5245]<=8'd232;
		data_a[5246]<=8'd231;
		data_a[5247]<=8'd230;
		data_a[5248]<=8'd228;
		data_a[5249]<=8'd227;
		data_a[5250]<=8'd254;
		data_a[5251]<=8'd196;
		data_a[5252]<=8'd187;
		data_a[5253]<=8'd173;
		data_a[5254]<=8'd208;
		data_a[5255]<=8'd191;
		data_a[5256]<=8'd201;
		data_a[5257]<=8'd202;
		data_a[5258]<=8'd203;
		data_a[5259]<=8'd210;
		data_a[5260]<=8'd215;
		data_a[5261]<=8'd215;
		data_a[5262]<=8'd213;
		data_a[5263]<=8'd214;
		data_a[5264]<=8'd208;
		data_a[5265]<=8'd209;
		data_a[5266]<=8'd210;
		data_a[5267]<=8'd210;
		data_a[5268]<=8'd210;
		data_a[5269]<=8'd208;
		data_a[5270]<=8'd210;
		data_a[5271]<=8'd209;
		data_a[5272]<=8'd204;
		data_a[5273]<=8'd203;
		data_a[5274]<=8'd206;
		data_a[5275]<=8'd200;
		data_a[5276]<=8'd135;
		data_a[5277]<=8'd194;
		data_a[5278]<=8'd183;
		data_a[5279]<=8'd168;
		data_a[5280]<=8'd121;
		data_a[5281]<=8'd90;
		data_a[5282]<=8'd86;
		data_a[5283]<=8'd109;
		data_a[5284]<=8'd105;
		data_a[5285]<=8'd97;
		data_a[5286]<=8'd78;
		data_a[5287]<=8'd90;
		data_a[5288]<=8'd80;
		data_a[5289]<=8'd83;
		data_a[5290]<=8'd74;
		data_a[5291]<=8'd73;
		data_a[5292]<=8'd77;
		data_a[5293]<=8'd73;
		data_a[5294]<=8'd71;
		data_a[5295]<=8'd79;
		data_a[5296]<=8'd83;
		data_a[5297]<=8'd89;
		data_a[5298]<=8'd92;
		data_a[5299]<=8'd106;
		data_a[5300]<=8'd104;
		data_a[5301]<=8'd119;
		data_a[5302]<=8'd120;
		data_a[5303]<=8'd119;
		data_a[5304]<=8'd115;
		data_a[5305]<=8'd109;
		data_a[5306]<=8'd102;
		data_a[5307]<=8'd108;
		data_a[5308]<=8'd119;
		data_a[5309]<=8'd113;
		data_a[5310]<=8'd122;
		data_a[5311]<=8'd133;
		data_a[5312]<=8'd113;
		data_a[5313]<=8'd114;
		data_a[5314]<=8'd141;
		data_a[5315]<=8'd221;
		data_a[5316]<=8'd218;
		data_a[5317]<=8'd213;
		data_a[5318]<=8'd209;
		data_a[5319]<=8'd215;
		data_a[5320]<=8'd217;
		data_a[5321]<=8'd216;
		data_a[5322]<=8'd213;
		data_a[5323]<=8'd212;
		data_a[5324]<=8'd212;
		data_a[5325]<=8'd208;
		data_a[5326]<=8'd218;
		data_a[5327]<=8'd182;
		data_a[5328]<=8'd89;
		data_a[5329]<=8'd101;
		data_a[5330]<=8'd96;
		data_a[5331]<=8'd85;
		data_a[5332]<=8'd79;
		data_a[5333]<=8'd74;
		data_a[5334]<=8'd75;
		data_a[5335]<=8'd66;
		data_a[5336]<=8'd71;
		data_a[5337]<=8'd74;
		data_a[5338]<=8'd86;
		data_a[5339]<=8'd92;
		data_a[5340]<=8'd102;
		data_a[5341]<=8'd110;
		data_a[5342]<=8'd120;
		data_a[5343]<=8'd130;
		data_a[5344]<=8'd138;
		data_a[5345]<=8'd149;
		data_a[5346]<=8'd160;
		data_a[5347]<=8'd167;
		data_a[5348]<=8'd170;
		data_a[5349]<=8'd170;
		data_a[5350]<=8'd171;
		data_a[5351]<=8'd172;
		data_a[5352]<=8'd171;
		data_a[5353]<=8'd172;
		data_a[5354]<=8'd176;
		data_a[5355]<=8'd178;
		data_a[5356]<=8'd181;
		data_a[5357]<=8'd183;
		data_a[5358]<=8'd182;
		data_a[5359]<=8'd180;
		data_a[5360]<=8'd179;
		data_a[5361]<=8'd180;
		data_a[5362]<=8'd180;
		data_a[5363]<=8'd183;
		data_a[5364]<=8'd182;
		data_a[5365]<=8'd174;
		data_a[5366]<=8'd171;
		data_a[5367]<=8'd160;
		data_a[5368]<=8'd145;
		data_a[5369]<=8'd119;
		data_a[5370]<=8'd112;
		data_a[5371]<=8'd111;
		data_a[5372]<=8'd128;
		data_a[5373]<=8'd141;
		data_a[5374]<=8'd206;
		data_a[5375]<=8'd216;
		data_a[5376]<=8'd218;
		data_a[5377]<=8'd217;
		data_a[5378]<=8'd218;
		data_a[5379]<=8'd218;
		data_a[5380]<=8'd222;
		data_a[5381]<=8'd221;
		data_a[5382]<=8'd226;
		data_a[5383]<=8'd225;
		data_a[5384]<=8'd228;
		data_a[5385]<=8'd227;
		data_a[5386]<=8'd228;
		data_a[5387]<=8'd227;
		data_a[5388]<=8'd228;
		data_a[5389]<=8'd229;
		data_a[5390]<=8'd230;
		data_a[5391]<=8'd229;
		data_a[5392]<=8'd230;
		data_a[5393]<=8'd231;
		data_a[5394]<=8'd230;
		data_a[5395]<=8'd230;
		data_a[5396]<=8'd230;
		data_a[5397]<=8'd229;
		data_a[5398]<=8'd227;
		data_a[5399]<=8'd226;
		data_a[5400]<=8'd251;
		data_a[5401]<=8'd201;
		data_a[5402]<=8'd203;
		data_a[5403]<=8'd164;
		data_a[5404]<=8'd204;
		data_a[5405]<=8'd186;
		data_a[5406]<=8'd205;
		data_a[5407]<=8'd207;
		data_a[5408]<=8'd212;
		data_a[5409]<=8'd212;
		data_a[5410]<=8'd215;
		data_a[5411]<=8'd208;
		data_a[5412]<=8'd209;
		data_a[5413]<=8'd214;
		data_a[5414]<=8'd215;
		data_a[5415]<=8'd211;
		data_a[5416]<=8'd209;
		data_a[5417]<=8'd209;
		data_a[5418]<=8'd208;
		data_a[5419]<=8'd206;
		data_a[5420]<=8'd208;
		data_a[5421]<=8'd208;
		data_a[5422]<=8'd203;
		data_a[5423]<=8'd202;
		data_a[5424]<=8'd203;
		data_a[5425]<=8'd201;
		data_a[5426]<=8'd189;
		data_a[5427]<=8'd189;
		data_a[5428]<=8'd182;
		data_a[5429]<=8'd159;
		data_a[5430]<=8'd136;
		data_a[5431]<=8'd105;
		data_a[5432]<=8'd89;
		data_a[5433]<=8'd98;
		data_a[5434]<=8'd106;
		data_a[5435]<=8'd103;
		data_a[5436]<=8'd82;
		data_a[5437]<=8'd86;
		data_a[5438]<=8'd83;
		data_a[5439]<=8'd81;
		data_a[5440]<=8'd77;
		data_a[5441]<=8'd71;
		data_a[5442]<=8'd74;
		data_a[5443]<=8'd72;
		data_a[5444]<=8'd76;
		data_a[5445]<=8'd84;
		data_a[5446]<=8'd84;
		data_a[5447]<=8'd84;
		data_a[5448]<=8'd95;
		data_a[5449]<=8'd94;
		data_a[5450]<=8'd96;
		data_a[5451]<=8'd109;
		data_a[5452]<=8'd110;
		data_a[5453]<=8'd107;
		data_a[5454]<=8'd115;
		data_a[5455]<=8'd108;
		data_a[5456]<=8'd100;
		data_a[5457]<=8'd105;
		data_a[5458]<=8'd100;
		data_a[5459]<=8'd117;
		data_a[5460]<=8'd98;
		data_a[5461]<=8'd110;
		data_a[5462]<=8'd103;
		data_a[5463]<=8'd110;
		data_a[5464]<=8'd142;
		data_a[5465]<=8'd187;
		data_a[5466]<=8'd207;
		data_a[5467]<=8'd214;
		data_a[5468]<=8'd215;
		data_a[5469]<=8'd208;
		data_a[5470]<=8'd218;
		data_a[5471]<=8'd214;
		data_a[5472]<=8'd212;
		data_a[5473]<=8'd216;
		data_a[5474]<=8'd208;
		data_a[5475]<=8'd210;
		data_a[5476]<=8'd217;
		data_a[5477]<=8'd138;
		data_a[5478]<=8'd111;
		data_a[5479]<=8'd90;
		data_a[5480]<=8'd91;
		data_a[5481]<=8'd85;
		data_a[5482]<=8'd75;
		data_a[5483]<=8'd71;
		data_a[5484]<=8'd70;
		data_a[5485]<=8'd75;
		data_a[5486]<=8'd69;
		data_a[5487]<=8'd84;
		data_a[5488]<=8'd95;
		data_a[5489]<=8'd101;
		data_a[5490]<=8'd112;
		data_a[5491]<=8'd119;
		data_a[5492]<=8'd129;
		data_a[5493]<=8'd140;
		data_a[5494]<=8'd146;
		data_a[5495]<=8'd153;
		data_a[5496]<=8'd165;
		data_a[5497]<=8'd170;
		data_a[5498]<=8'd172;
		data_a[5499]<=8'd172;
		data_a[5500]<=8'd175;
		data_a[5501]<=8'd176;
		data_a[5502]<=8'd175;
		data_a[5503]<=8'd174;
		data_a[5504]<=8'd173;
		data_a[5505]<=8'd179;
		data_a[5506]<=8'd184;
		data_a[5507]<=8'd184;
		data_a[5508]<=8'd182;
		data_a[5509]<=8'd182;
		data_a[5510]<=8'd179;
		data_a[5511]<=8'd177;
		data_a[5512]<=8'd176;
		data_a[5513]<=8'd179;
		data_a[5514]<=8'd187;
		data_a[5515]<=8'd178;
		data_a[5516]<=8'd177;
		data_a[5517]<=8'd170;
		data_a[5518]<=8'd151;
		data_a[5519]<=8'd124;
		data_a[5520]<=8'd109;
		data_a[5521]<=8'd111;
		data_a[5522]<=8'd126;
		data_a[5523]<=8'd147;
		data_a[5524]<=8'd186;
		data_a[5525]<=8'd214;
		data_a[5526]<=8'd217;
		data_a[5527]<=8'd219;
		data_a[5528]<=8'd218;
		data_a[5529]<=8'd218;
		data_a[5530]<=8'd221;
		data_a[5531]<=8'd220;
		data_a[5532]<=8'd225;
		data_a[5533]<=8'd223;
		data_a[5534]<=8'd226;
		data_a[5535]<=8'd226;
		data_a[5536]<=8'd227;
		data_a[5537]<=8'd227;
		data_a[5538]<=8'd228;
		data_a[5539]<=8'd229;
		data_a[5540]<=8'd230;
		data_a[5541]<=8'd229;
		data_a[5542]<=8'd229;
		data_a[5543]<=8'd229;
		data_a[5544]<=8'd229;
		data_a[5545]<=8'd229;
		data_a[5546]<=8'd230;
		data_a[5547]<=8'd230;
		data_a[5548]<=8'd229;
		data_a[5549]<=8'd227;
		data_a[5550]<=8'd254;
		data_a[5551]<=8'd202;
		data_a[5552]<=8'd202;
		data_a[5553]<=8'd192;
		data_a[5554]<=8'd209;
		data_a[5555]<=8'd217;
		data_a[5556]<=8'd214;
		data_a[5557]<=8'd215;
		data_a[5558]<=8'd211;
		data_a[5559]<=8'd215;
		data_a[5560]<=8'd209;
		data_a[5561]<=8'd212;
		data_a[5562]<=8'd213;
		data_a[5563]<=8'd212;
		data_a[5564]<=8'd209;
		data_a[5565]<=8'd212;
		data_a[5566]<=8'd211;
		data_a[5567]<=8'd209;
		data_a[5568]<=8'd207;
		data_a[5569]<=8'd207;
		data_a[5570]<=8'd207;
		data_a[5571]<=8'd207;
		data_a[5572]<=8'd205;
		data_a[5573]<=8'd201;
		data_a[5574]<=8'd193;
		data_a[5575]<=8'd176;
		data_a[5576]<=8'd137;
		data_a[5577]<=8'd140;
		data_a[5578]<=8'd137;
		data_a[5579]<=8'd166;
		data_a[5580]<=8'd139;
		data_a[5581]<=8'd133;
		data_a[5582]<=8'd84;
		data_a[5583]<=8'd103;
		data_a[5584]<=8'd90;
		data_a[5585]<=8'd87;
		data_a[5586]<=8'd85;
		data_a[5587]<=8'd78;
		data_a[5588]<=8'd84;
		data_a[5589]<=8'd83;
		data_a[5590]<=8'd73;
		data_a[5591]<=8'd69;
		data_a[5592]<=8'd74;
		data_a[5593]<=8'd77;
		data_a[5594]<=8'd82;
		data_a[5595]<=8'd81;
		data_a[5596]<=8'd79;
		data_a[5597]<=8'd75;
		data_a[5598]<=8'd103;
		data_a[5599]<=8'd89;
		data_a[5600]<=8'd97;
		data_a[5601]<=8'd100;
		data_a[5602]<=8'd99;
		data_a[5603]<=8'd101;
		data_a[5604]<=8'd109;
		data_a[5605]<=8'd108;
		data_a[5606]<=8'd95;
		data_a[5607]<=8'd109;
		data_a[5608]<=8'd94;
		data_a[5609]<=8'd110;
		data_a[5610]<=8'd107;
		data_a[5611]<=8'd93;
		data_a[5612]<=8'd96;
		data_a[5613]<=8'd106;
		data_a[5614]<=8'd127;
		data_a[5615]<=8'd146;
		data_a[5616]<=8'd221;
		data_a[5617]<=8'd211;
		data_a[5618]<=8'd215;
		data_a[5619]<=8'd213;
		data_a[5620]<=8'd214;
		data_a[5621]<=8'd215;
		data_a[5622]<=8'd212;
		data_a[5623]<=8'd213;
		data_a[5624]<=8'd209;
		data_a[5625]<=8'd213;
		data_a[5626]<=8'd209;
		data_a[5627]<=8'd86;
		data_a[5628]<=8'd99;
		data_a[5629]<=8'd98;
		data_a[5630]<=8'd88;
		data_a[5631]<=8'd75;
		data_a[5632]<=8'd74;
		data_a[5633]<=8'd64;
		data_a[5634]<=8'd62;
		data_a[5635]<=8'd72;
		data_a[5636]<=8'd79;
		data_a[5637]<=8'd94;
		data_a[5638]<=8'd102;
		data_a[5639]<=8'd110;
		data_a[5640]<=8'd121;
		data_a[5641]<=8'd126;
		data_a[5642]<=8'd137;
		data_a[5643]<=8'd148;
		data_a[5644]<=8'd151;
		data_a[5645]<=8'd155;
		data_a[5646]<=8'd164;
		data_a[5647]<=8'd170;
		data_a[5648]<=8'd173;
		data_a[5649]<=8'd173;
		data_a[5650]<=8'd174;
		data_a[5651]<=8'd174;
		data_a[5652]<=8'd174;
		data_a[5653]<=8'd175;
		data_a[5654]<=8'd172;
		data_a[5655]<=8'd178;
		data_a[5656]<=8'd181;
		data_a[5657]<=8'd178;
		data_a[5658]<=8'd177;
		data_a[5659]<=8'd179;
		data_a[5660]<=8'd180;
		data_a[5661]<=8'd178;
		data_a[5662]<=8'd185;
		data_a[5663]<=8'd174;
		data_a[5664]<=8'd184;
		data_a[5665]<=8'd181;
		data_a[5666]<=8'd177;
		data_a[5667]<=8'd175;
		data_a[5668]<=8'd163;
		data_a[5669]<=8'd134;
		data_a[5670]<=8'd113;
		data_a[5671]<=8'd117;
		data_a[5672]<=8'd125;
		data_a[5673]<=8'd132;
		data_a[5674]<=8'd201;
		data_a[5675]<=8'd217;
		data_a[5676]<=8'd210;
		data_a[5677]<=8'd218;
		data_a[5678]<=8'd218;
		data_a[5679]<=8'd218;
		data_a[5680]<=8'd220;
		data_a[5681]<=8'd220;
		data_a[5682]<=8'd222;
		data_a[5683]<=8'd221;
		data_a[5684]<=8'd223;
		data_a[5685]<=8'd224;
		data_a[5686]<=8'd225;
		data_a[5687]<=8'd226;
		data_a[5688]<=8'd227;
		data_a[5689]<=8'd228;
		data_a[5690]<=8'd228;
		data_a[5691]<=8'd228;
		data_a[5692]<=8'd228;
		data_a[5693]<=8'd228;
		data_a[5694]<=8'd229;
		data_a[5695]<=8'd230;
		data_a[5696]<=8'd231;
		data_a[5697]<=8'd231;
		data_a[5698]<=8'd230;
		data_a[5699]<=8'd229;
		data_a[5700]<=8'd255;
		data_a[5701]<=8'd206;
		data_a[5702]<=8'd214;
		data_a[5703]<=8'd214;
		data_a[5704]<=8'd214;
		data_a[5705]<=8'd218;
		data_a[5706]<=8'd212;
		data_a[5707]<=8'd213;
		data_a[5708]<=8'd212;
		data_a[5709]<=8'd207;
		data_a[5710]<=8'd211;
		data_a[5711]<=8'd211;
		data_a[5712]<=8'd210;
		data_a[5713]<=8'd212;
		data_a[5714]<=8'd207;
		data_a[5715]<=8'd218;
		data_a[5716]<=8'd211;
		data_a[5717]<=8'd210;
		data_a[5718]<=8'd207;
		data_a[5719]<=8'd208;
		data_a[5720]<=8'd204;
		data_a[5721]<=8'd199;
		data_a[5722]<=8'd198;
		data_a[5723]<=8'd188;
		data_a[5724]<=8'd184;
		data_a[5725]<=8'd185;
		data_a[5726]<=8'd168;
		data_a[5727]<=8'd191;
		data_a[5728]<=8'd179;
		data_a[5729]<=8'd175;
		data_a[5730]<=8'd132;
		data_a[5731]<=8'd123;
		data_a[5732]<=8'd99;
		data_a[5733]<=8'd112;
		data_a[5734]<=8'd98;
		data_a[5735]<=8'd82;
		data_a[5736]<=8'd90;
		data_a[5737]<=8'd92;
		data_a[5738]<=8'd85;
		data_a[5739]<=8'd92;
		data_a[5740]<=8'd72;
		data_a[5741]<=8'd71;
		data_a[5742]<=8'd74;
		data_a[5743]<=8'd73;
		data_a[5744]<=8'd71;
		data_a[5745]<=8'd67;
		data_a[5746]<=8'd77;
		data_a[5747]<=8'd82;
		data_a[5748]<=8'd93;
		data_a[5749]<=8'd89;
		data_a[5750]<=8'd97;
		data_a[5751]<=8'd96;
		data_a[5752]<=8'd92;
		data_a[5753]<=8'd95;
		data_a[5754]<=8'd102;
		data_a[5755]<=8'd104;
		data_a[5756]<=8'd94;
		data_a[5757]<=8'd92;
		data_a[5758]<=8'd92;
		data_a[5759]<=8'd99;
		data_a[5760]<=8'd101;
		data_a[5761]<=8'd90;
		data_a[5762]<=8'd97;
		data_a[5763]<=8'd98;
		data_a[5764]<=8'd116;
		data_a[5765]<=8'd132;
		data_a[5766]<=8'd223;
		data_a[5767]<=8'd212;
		data_a[5768]<=8'd214;
		data_a[5769]<=8'd220;
		data_a[5770]<=8'd211;
		data_a[5771]<=8'd213;
		data_a[5772]<=8'd215;
		data_a[5773]<=8'd211;
		data_a[5774]<=8'd211;
		data_a[5775]<=8'd205;
		data_a[5776]<=8'd213;
		data_a[5777]<=8'd100;
		data_a[5778]<=8'd88;
		data_a[5779]<=8'd80;
		data_a[5780]<=8'd79;
		data_a[5781]<=8'd69;
		data_a[5782]<=8'd72;
		data_a[5783]<=8'd70;
		data_a[5784]<=8'd69;
		data_a[5785]<=8'd80;
		data_a[5786]<=8'd93;
		data_a[5787]<=8'd100;
		data_a[5788]<=8'd111;
		data_a[5789]<=8'd121;
		data_a[5790]<=8'd131;
		data_a[5791]<=8'd134;
		data_a[5792]<=8'd143;
		data_a[5793]<=8'd154;
		data_a[5794]<=8'd156;
		data_a[5795]<=8'd158;
		data_a[5796]<=8'd164;
		data_a[5797]<=8'd170;
		data_a[5798]<=8'd171;
		data_a[5799]<=8'd171;
		data_a[5800]<=8'd172;
		data_a[5801]<=8'd172;
		data_a[5802]<=8'd172;
		data_a[5803]<=8'd173;
		data_a[5804]<=8'd173;
		data_a[5805]<=8'd175;
		data_a[5806]<=8'd176;
		data_a[5807]<=8'd173;
		data_a[5808]<=8'd172;
		data_a[5809]<=8'd176;
		data_a[5810]<=8'd179;
		data_a[5811]<=8'd180;
		data_a[5812]<=8'd181;
		data_a[5813]<=8'd177;
		data_a[5814]<=8'd182;
		data_a[5815]<=8'd186;
		data_a[5816]<=8'd183;
		data_a[5817]<=8'd180;
		data_a[5818]<=8'd172;
		data_a[5819]<=8'd143;
		data_a[5820]<=8'd114;
		data_a[5821]<=8'd123;
		data_a[5822]<=8'd122;
		data_a[5823]<=8'd131;
		data_a[5824]<=8'd159;
		data_a[5825]<=8'd215;
		data_a[5826]<=8'd216;
		data_a[5827]<=8'd217;
		data_a[5828]<=8'd217;
		data_a[5829]<=8'd218;
		data_a[5830]<=8'd219;
		data_a[5831]<=8'd221;
		data_a[5832]<=8'd220;
		data_a[5833]<=8'd220;
		data_a[5834]<=8'd221;
		data_a[5835]<=8'd223;
		data_a[5836]<=8'd223;
		data_a[5837]<=8'd224;
		data_a[5838]<=8'd225;
		data_a[5839]<=8'd226;
		data_a[5840]<=8'd226;
		data_a[5841]<=8'd227;
		data_a[5842]<=8'd227;
		data_a[5843]<=8'd227;
		data_a[5844]<=8'd229;
		data_a[5845]<=8'd230;
		data_a[5846]<=8'd231;
		data_a[5847]<=8'd231;
		data_a[5848]<=8'd230;
		data_a[5849]<=8'd230;
		data_a[5850]<=8'd255;
		data_a[5851]<=8'd212;
		data_a[5852]<=8'd216;
		data_a[5853]<=8'd218;
		data_a[5854]<=8'd211;
		data_a[5855]<=8'd212;
		data_a[5856]<=8'd212;
		data_a[5857]<=8'd213;
		data_a[5858]<=8'd212;
		data_a[5859]<=8'd212;
		data_a[5860]<=8'd209;
		data_a[5861]<=8'd213;
		data_a[5862]<=8'd206;
		data_a[5863]<=8'd209;
		data_a[5864]<=8'd213;
		data_a[5865]<=8'd209;
		data_a[5866]<=8'd208;
		data_a[5867]<=8'd208;
		data_a[5868]<=8'd205;
		data_a[5869]<=8'd209;
		data_a[5870]<=8'd200;
		data_a[5871]<=8'd190;
		data_a[5872]<=8'd186;
		data_a[5873]<=8'd170;
		data_a[5874]<=8'd163;
		data_a[5875]<=8'd149;
		data_a[5876]<=8'd158;
		data_a[5877]<=8'd118;
		data_a[5878]<=8'd159;
		data_a[5879]<=8'd152;
		data_a[5880]<=8'd129;
		data_a[5881]<=8'd118;
		data_a[5882]<=8'd96;
		data_a[5883]<=8'd102;
		data_a[5884]<=8'd88;
		data_a[5885]<=8'd89;
		data_a[5886]<=8'd83;
		data_a[5887]<=8'd83;
		data_a[5888]<=8'd91;
		data_a[5889]<=8'd72;
		data_a[5890]<=8'd69;
		data_a[5891]<=8'd70;
		data_a[5892]<=8'd72;
		data_a[5893]<=8'd71;
		data_a[5894]<=8'd67;
		data_a[5895]<=8'd59;
		data_a[5896]<=8'd75;
		data_a[5897]<=8'd83;
		data_a[5898]<=8'd87;
		data_a[5899]<=8'd86;
		data_a[5900]<=8'd77;
		data_a[5901]<=8'd92;
		data_a[5902]<=8'd104;
		data_a[5903]<=8'd111;
		data_a[5904]<=8'd109;
		data_a[5905]<=8'd93;
		data_a[5906]<=8'd100;
		data_a[5907]<=8'd91;
		data_a[5908]<=8'd93;
		data_a[5909]<=8'd101;
		data_a[5910]<=8'd94;
		data_a[5911]<=8'd101;
		data_a[5912]<=8'd88;
		data_a[5913]<=8'd114;
		data_a[5914]<=8'd122;
		data_a[5915]<=8'd140;
		data_a[5916]<=8'd189;
		data_a[5917]<=8'd210;
		data_a[5918]<=8'd214;
		data_a[5919]<=8'd213;
		data_a[5920]<=8'd214;
		data_a[5921]<=8'd210;
		data_a[5922]<=8'd207;
		data_a[5923]<=8'd210;
		data_a[5924]<=8'd213;
		data_a[5925]<=8'd208;
		data_a[5926]<=8'd194;
		data_a[5927]<=8'd84;
		data_a[5928]<=8'd87;
		data_a[5929]<=8'd80;
		data_a[5930]<=8'd75;
		data_a[5931]<=8'd72;
		data_a[5932]<=8'd61;
		data_a[5933]<=8'd71;
		data_a[5934]<=8'd72;
		data_a[5935]<=8'd90;
		data_a[5936]<=8'd100;
		data_a[5937]<=8'd109;
		data_a[5938]<=8'd119;
		data_a[5939]<=8'd130;
		data_a[5940]<=8'd139;
		data_a[5941]<=8'd141;
		data_a[5942]<=8'd148;
		data_a[5943]<=8'd159;
		data_a[5944]<=8'd160;
		data_a[5945]<=8'd162;
		data_a[5946]<=8'd168;
		data_a[5947]<=8'd171;
		data_a[5948]<=8'd170;
		data_a[5949]<=8'd169;
		data_a[5950]<=8'd172;
		data_a[5951]<=8'd174;
		data_a[5952]<=8'd172;
		data_a[5953]<=8'd171;
		data_a[5954]<=8'd169;
		data_a[5955]<=8'd172;
		data_a[5956]<=8'd175;
		data_a[5957]<=8'd176;
		data_a[5958]<=8'd176;
		data_a[5959]<=8'd176;
		data_a[5960]<=8'd177;
		data_a[5961]<=8'd178;
		data_a[5962]<=8'd174;
		data_a[5963]<=8'd187;
		data_a[5964]<=8'd181;
		data_a[5965]<=8'd182;
		data_a[5966]<=8'd185;
		data_a[5967]<=8'd183;
		data_a[5968]<=8'd177;
		data_a[5969]<=8'd154;
		data_a[5970]<=8'd124;
		data_a[5971]<=8'd119;
		data_a[5972]<=8'd113;
		data_a[5973]<=8'd135;
		data_a[5974]<=8'd143;
		data_a[5975]<=8'd214;
		data_a[5976]<=8'd217;
		data_a[5977]<=8'd217;
		data_a[5978]<=8'd217;
		data_a[5979]<=8'd218;
		data_a[5980]<=8'd218;
		data_a[5981]<=8'd222;
		data_a[5982]<=8'd218;
		data_a[5983]<=8'd220;
		data_a[5984]<=8'd219;
		data_a[5985]<=8'd222;
		data_a[5986]<=8'd223;
		data_a[5987]<=8'd224;
		data_a[5988]<=8'd225;
		data_a[5989]<=8'd225;
		data_a[5990]<=8'd226;
		data_a[5991]<=8'd227;
		data_a[5992]<=8'd228;
		data_a[5993]<=8'd229;
		data_a[5994]<=8'd228;
		data_a[5995]<=8'd229;
		data_a[5996]<=8'd229;
		data_a[5997]<=8'd229;
		data_a[5998]<=8'd228;
		data_a[5999]<=8'd229;
		data_a[6000]<=8'd255;
		data_a[6001]<=8'd212;
		data_a[6002]<=8'd214;
		data_a[6003]<=8'd211;
		data_a[6004]<=8'd212;
		data_a[6005]<=8'd214;
		data_a[6006]<=8'd214;
		data_a[6007]<=8'd207;
		data_a[6008]<=8'd209;
		data_a[6009]<=8'd211;
		data_a[6010]<=8'd212;
		data_a[6011]<=8'd211;
		data_a[6012]<=8'd210;
		data_a[6013]<=8'd210;
		data_a[6014]<=8'd210;
		data_a[6015]<=8'd209;
		data_a[6016]<=8'd211;
		data_a[6017]<=8'd208;
		data_a[6018]<=8'd202;
		data_a[6019]<=8'd196;
		data_a[6020]<=8'd196;
		data_a[6021]<=8'd195;
		data_a[6022]<=8'd206;
		data_a[6023]<=8'd171;
		data_a[6024]<=8'd159;
		data_a[6025]<=8'd123;
		data_a[6026]<=8'd99;
		data_a[6027]<=8'd127;
		data_a[6028]<=8'd116;
		data_a[6029]<=8'd118;
		data_a[6030]<=8'd107;
		data_a[6031]<=8'd105;
		data_a[6032]<=8'd92;
		data_a[6033]<=8'd94;
		data_a[6034]<=8'd80;
		data_a[6035]<=8'd77;
		data_a[6036]<=8'd79;
		data_a[6037]<=8'd80;
		data_a[6038]<=8'd81;
		data_a[6039]<=8'd81;
		data_a[6040]<=8'd70;
		data_a[6041]<=8'd69;
		data_a[6042]<=8'd71;
		data_a[6043]<=8'd73;
		data_a[6044]<=8'd70;
		data_a[6045]<=8'd76;
		data_a[6046]<=8'd73;
		data_a[6047]<=8'd80;
		data_a[6048]<=8'd83;
		data_a[6049]<=8'd76;
		data_a[6050]<=8'd77;
		data_a[6051]<=8'd94;
		data_a[6052]<=8'd100;
		data_a[6053]<=8'd97;
		data_a[6054]<=8'd99;
		data_a[6055]<=8'd97;
		data_a[6056]<=8'd95;
		data_a[6057]<=8'd96;
		data_a[6058]<=8'd99;
		data_a[6059]<=8'd92;
		data_a[6060]<=8'd92;
		data_a[6061]<=8'd94;
		data_a[6062]<=8'd85;
		data_a[6063]<=8'd119;
		data_a[6064]<=8'd97;
		data_a[6065]<=8'd166;
		data_a[6066]<=8'd189;
		data_a[6067]<=8'd204;
		data_a[6068]<=8'd211;
		data_a[6069]<=8'd207;
		data_a[6070]<=8'd213;
		data_a[6071]<=8'd212;
		data_a[6072]<=8'd211;
		data_a[6073]<=8'd209;
		data_a[6074]<=8'd212;
		data_a[6075]<=8'd207;
		data_a[6076]<=8'd204;
		data_a[6077]<=8'd75;
		data_a[6078]<=8'd81;
		data_a[6079]<=8'd77;
		data_a[6080]<=8'd75;
		data_a[6081]<=8'd66;
		data_a[6082]<=8'd65;
		data_a[6083]<=8'd65;
		data_a[6084]<=8'd72;
		data_a[6085]<=8'd99;
		data_a[6086]<=8'd109;
		data_a[6087]<=8'd121;
		data_a[6088]<=8'd131;
		data_a[6089]<=8'd138;
		data_a[6090]<=8'd142;
		data_a[6091]<=8'd151;
		data_a[6092]<=8'd157;
		data_a[6093]<=8'd158;
		data_a[6094]<=8'd165;
		data_a[6095]<=8'd165;
		data_a[6096]<=8'd164;
		data_a[6097]<=8'd164;
		data_a[6098]<=8'd166;
		data_a[6099]<=8'd169;
		data_a[6100]<=8'd170;
		data_a[6101]<=8'd173;
		data_a[6102]<=8'd173;
		data_a[6103]<=8'd170;
		data_a[6104]<=8'd173;
		data_a[6105]<=8'd169;
		data_a[6106]<=8'd171;
		data_a[6107]<=8'd171;
		data_a[6108]<=8'd178;
		data_a[6109]<=8'd176;
		data_a[6110]<=8'd179;
		data_a[6111]<=8'd179;
		data_a[6112]<=8'd180;
		data_a[6113]<=8'd178;
		data_a[6114]<=8'd181;
		data_a[6115]<=8'd182;
		data_a[6116]<=8'd183;
		data_a[6117]<=8'd188;
		data_a[6118]<=8'd181;
		data_a[6119]<=8'd162;
		data_a[6120]<=8'd128;
		data_a[6121]<=8'd116;
		data_a[6122]<=8'd118;
		data_a[6123]<=8'd131;
		data_a[6124]<=8'd125;
		data_a[6125]<=8'd196;
		data_a[6126]<=8'd219;
		data_a[6127]<=8'd214;
		data_a[6128]<=8'd213;
		data_a[6129]<=8'd218;
		data_a[6130]<=8'd220;
		data_a[6131]<=8'd219;
		data_a[6132]<=8'd219;
		data_a[6133]<=8'd223;
		data_a[6134]<=8'd224;
		data_a[6135]<=8'd223;
		data_a[6136]<=8'd223;
		data_a[6137]<=8'd224;
		data_a[6138]<=8'd225;
		data_a[6139]<=8'd226;
		data_a[6140]<=8'd226;
		data_a[6141]<=8'd227;
		data_a[6142]<=8'd229;
		data_a[6143]<=8'd231;
		data_a[6144]<=8'd229;
		data_a[6145]<=8'd230;
		data_a[6146]<=8'd230;
		data_a[6147]<=8'd230;
		data_a[6148]<=8'd230;
		data_a[6149]<=8'd230;
		data_a[6150]<=8'd255;
		data_a[6151]<=8'd215;
		data_a[6152]<=8'd211;
		data_a[6153]<=8'd210;
		data_a[6154]<=8'd215;
		data_a[6155]<=8'd208;
		data_a[6156]<=8'd206;
		data_a[6157]<=8'd215;
		data_a[6158]<=8'd210;
		data_a[6159]<=8'd212;
		data_a[6160]<=8'd212;
		data_a[6161]<=8'd211;
		data_a[6162]<=8'd210;
		data_a[6163]<=8'd209;
		data_a[6164]<=8'd209;
		data_a[6165]<=8'd208;
		data_a[6166]<=8'd206;
		data_a[6167]<=8'd206;
		data_a[6168]<=8'd190;
		data_a[6169]<=8'd202;
		data_a[6170]<=8'd192;
		data_a[6171]<=8'd188;
		data_a[6172]<=8'd178;
		data_a[6173]<=8'd162;
		data_a[6174]<=8'd160;
		data_a[6175]<=8'd113;
		data_a[6176]<=8'd112;
		data_a[6177]<=8'd102;
		data_a[6178]<=8'd87;
		data_a[6179]<=8'd94;
		data_a[6180]<=8'd90;
		data_a[6181]<=8'd88;
		data_a[6182]<=8'd87;
		data_a[6183]<=8'd83;
		data_a[6184]<=8'd82;
		data_a[6185]<=8'd78;
		data_a[6186]<=8'd81;
		data_a[6187]<=8'd76;
		data_a[6188]<=8'd75;
		data_a[6189]<=8'd67;
		data_a[6190]<=8'd68;
		data_a[6191]<=8'd67;
		data_a[6192]<=8'd70;
		data_a[6193]<=8'd68;
		data_a[6194]<=8'd69;
		data_a[6195]<=8'd73;
		data_a[6196]<=8'd71;
		data_a[6197]<=8'd73;
		data_a[6198]<=8'd75;
		data_a[6199]<=8'd72;
		data_a[6200]<=8'd75;
		data_a[6201]<=8'd88;
		data_a[6202]<=8'd93;
		data_a[6203]<=8'd94;
		data_a[6204]<=8'd100;
		data_a[6205]<=8'd98;
		data_a[6206]<=8'd97;
		data_a[6207]<=8'd91;
		data_a[6208]<=8'd94;
		data_a[6209]<=8'd94;
		data_a[6210]<=8'd94;
		data_a[6211]<=8'd92;
		data_a[6212]<=8'd85;
		data_a[6213]<=8'd85;
		data_a[6214]<=8'd96;
		data_a[6215]<=8'd182;
		data_a[6216]<=8'd179;
		data_a[6217]<=8'd204;
		data_a[6218]<=8'd210;
		data_a[6219]<=8'd212;
		data_a[6220]<=8'd210;
		data_a[6221]<=8'd211;
		data_a[6222]<=8'd212;
		data_a[6223]<=8'd212;
		data_a[6224]<=8'd206;
		data_a[6225]<=8'd213;
		data_a[6226]<=8'd196;
		data_a[6227]<=8'd93;
		data_a[6228]<=8'd81;
		data_a[6229]<=8'd76;
		data_a[6230]<=8'd76;
		data_a[6231]<=8'd66;
		data_a[6232]<=8'd62;
		data_a[6233]<=8'd66;
		data_a[6234]<=8'd83;
		data_a[6235]<=8'd104;
		data_a[6236]<=8'd115;
		data_a[6237]<=8'd129;
		data_a[6238]<=8'd139;
		data_a[6239]<=8'd144;
		data_a[6240]<=8'd149;
		data_a[6241]<=8'd156;
		data_a[6242]<=8'd160;
		data_a[6243]<=8'd162;
		data_a[6244]<=8'd166;
		data_a[6245]<=8'd166;
		data_a[6246]<=8'd163;
		data_a[6247]<=8'd163;
		data_a[6248]<=8'd165;
		data_a[6249]<=8'd167;
		data_a[6250]<=8'd168;
		data_a[6251]<=8'd171;
		data_a[6252]<=8'd172;
		data_a[6253]<=8'd169;
		data_a[6254]<=8'd163;
		data_a[6255]<=8'd165;
		data_a[6256]<=8'd172;
		data_a[6257]<=8'd174;
		data_a[6258]<=8'd179;
		data_a[6259]<=8'd177;
		data_a[6260]<=8'd179;
		data_a[6261]<=8'd179;
		data_a[6262]<=8'd180;
		data_a[6263]<=8'd178;
		data_a[6264]<=8'd180;
		data_a[6265]<=8'd180;
		data_a[6266]<=8'd180;
		data_a[6267]<=8'd186;
		data_a[6268]<=8'd182;
		data_a[6269]<=8'd167;
		data_a[6270]<=8'd132;
		data_a[6271]<=8'd121;
		data_a[6272]<=8'd116;
		data_a[6273]<=8'd122;
		data_a[6274]<=8'd133;
		data_a[6275]<=8'd149;
		data_a[6276]<=8'd212;
		data_a[6277]<=8'd214;
		data_a[6278]<=8'd214;
		data_a[6279]<=8'd218;
		data_a[6280]<=8'd221;
		data_a[6281]<=8'd220;
		data_a[6282]<=8'd220;
		data_a[6283]<=8'd223;
		data_a[6284]<=8'd224;
		data_a[6285]<=8'd222;
		data_a[6286]<=8'd225;
		data_a[6287]<=8'd223;
		data_a[6288]<=8'd221;
		data_a[6289]<=8'd221;
		data_a[6290]<=8'd224;
		data_a[6291]<=8'd228;
		data_a[6292]<=8'd230;
		data_a[6293]<=8'd230;
		data_a[6294]<=8'd230;
		data_a[6295]<=8'd231;
		data_a[6296]<=8'd230;
		data_a[6297]<=8'd229;
		data_a[6298]<=8'd230;
		data_a[6299]<=8'd231;
		data_a[6300]<=8'd254;
		data_a[6301]<=8'd210;
		data_a[6302]<=8'd210;
		data_a[6303]<=8'd210;
		data_a[6304]<=8'd210;
		data_a[6305]<=8'd212;
		data_a[6306]<=8'd212;
		data_a[6307]<=8'd209;
		data_a[6308]<=8'd210;
		data_a[6309]<=8'd212;
		data_a[6310]<=8'd212;
		data_a[6311]<=8'd210;
		data_a[6312]<=8'd209;
		data_a[6313]<=8'd209;
		data_a[6314]<=8'd208;
		data_a[6315]<=8'd208;
		data_a[6316]<=8'd211;
		data_a[6317]<=8'd212;
		data_a[6318]<=8'd184;
		data_a[6319]<=8'd213;
		data_a[6320]<=8'd189;
		data_a[6321]<=8'd176;
		data_a[6322]<=8'd146;
		data_a[6323]<=8'd143;
		data_a[6324]<=8'd120;
		data_a[6325]<=8'd98;
		data_a[6326]<=8'd113;
		data_a[6327]<=8'd128;
		data_a[6328]<=8'd85;
		data_a[6329]<=8'd85;
		data_a[6330]<=8'd87;
		data_a[6331]<=8'd80;
		data_a[6332]<=8'd81;
		data_a[6333]<=8'd75;
		data_a[6334]<=8'd73;
		data_a[6335]<=8'd77;
		data_a[6336]<=8'd68;
		data_a[6337]<=8'd75;
		data_a[6338]<=8'd71;
		data_a[6339]<=8'd67;
		data_a[6340]<=8'd67;
		data_a[6341]<=8'd69;
		data_a[6342]<=8'd68;
		data_a[6343]<=8'd70;
		data_a[6344]<=8'd67;
		data_a[6345]<=8'd75;
		data_a[6346]<=8'd71;
		data_a[6347]<=8'd72;
		data_a[6348]<=8'd75;
		data_a[6349]<=8'd78;
		data_a[6350]<=8'd80;
		data_a[6351]<=8'd85;
		data_a[6352]<=8'd85;
		data_a[6353]<=8'd87;
		data_a[6354]<=8'd93;
		data_a[6355]<=8'd93;
		data_a[6356]<=8'd93;
		data_a[6357]<=8'd91;
		data_a[6358]<=8'd92;
		data_a[6359]<=8'd97;
		data_a[6360]<=8'd101;
		data_a[6361]<=8'd98;
		data_a[6362]<=8'd103;
		data_a[6363]<=8'd92;
		data_a[6364]<=8'd96;
		data_a[6365]<=8'd140;
		data_a[6366]<=8'd173;
		data_a[6367]<=8'd202;
		data_a[6368]<=8'd208;
		data_a[6369]<=8'd212;
		data_a[6370]<=8'd207;
		data_a[6371]<=8'd210;
		data_a[6372]<=8'd204;
		data_a[6373]<=8'd218;
		data_a[6374]<=8'd211;
		data_a[6375]<=8'd208;
		data_a[6376]<=8'd206;
		data_a[6377]<=8'd83;
		data_a[6378]<=8'd84;
		data_a[6379]<=8'd79;
		data_a[6380]<=8'd73;
		data_a[6381]<=8'd66;
		data_a[6382]<=8'd61;
		data_a[6383]<=8'd73;
		data_a[6384]<=8'd96;
		data_a[6385]<=8'd111;
		data_a[6386]<=8'd123;
		data_a[6387]<=8'd139;
		data_a[6388]<=8'd144;
		data_a[6389]<=8'd147;
		data_a[6390]<=8'd154;
		data_a[6391]<=8'd158;
		data_a[6392]<=8'd162;
		data_a[6393]<=8'd165;
		data_a[6394]<=8'd164;
		data_a[6395]<=8'd166;
		data_a[6396]<=8'd171;
		data_a[6397]<=8'd170;
		data_a[6398]<=8'd172;
		data_a[6399]<=8'd172;
		data_a[6400]<=8'd171;
		data_a[6401]<=8'd171;
		data_a[6402]<=8'd169;
		data_a[6403]<=8'd166;
		data_a[6404]<=8'd151;
		data_a[6405]<=8'd159;
		data_a[6406]<=8'd171;
		data_a[6407]<=8'd175;
		data_a[6408]<=8'd180;
		data_a[6409]<=8'd179;
		data_a[6410]<=8'd181;
		data_a[6411]<=8'd181;
		data_a[6412]<=8'd179;
		data_a[6413]<=8'd179;
		data_a[6414]<=8'd181;
		data_a[6415]<=8'd180;
		data_a[6416]<=8'd180;
		data_a[6417]<=8'd185;
		data_a[6418]<=8'd183;
		data_a[6419]<=8'd172;
		data_a[6420]<=8'd143;
		data_a[6421]<=8'd119;
		data_a[6422]<=8'd120;
		data_a[6423]<=8'd116;
		data_a[6424]<=8'd124;
		data_a[6425]<=8'd140;
		data_a[6426]<=8'd195;
		data_a[6427]<=8'd209;
		data_a[6428]<=8'd215;
		data_a[6429]<=8'd218;
		data_a[6430]<=8'd220;
		data_a[6431]<=8'd220;
		data_a[6432]<=8'd220;
		data_a[6433]<=8'd222;
		data_a[6434]<=8'd223;
		data_a[6435]<=8'd221;
		data_a[6436]<=8'd224;
		data_a[6437]<=8'd223;
		data_a[6438]<=8'd222;
		data_a[6439]<=8'd223;
		data_a[6440]<=8'd226;
		data_a[6441]<=8'd228;
		data_a[6442]<=8'd228;
		data_a[6443]<=8'd227;
		data_a[6444]<=8'd227;
		data_a[6445]<=8'd229;
		data_a[6446]<=8'd230;
		data_a[6447]<=8'd231;
		data_a[6448]<=8'd232;
		data_a[6449]<=8'd232;
		data_a[6450]<=8'd255;
		data_a[6451]<=8'd208;
		data_a[6452]<=8'd211;
		data_a[6453]<=8'd214;
		data_a[6454]<=8'd208;
		data_a[6455]<=8'd211;
		data_a[6456]<=8'd213;
		data_a[6457]<=8'd210;
		data_a[6458]<=8'd210;
		data_a[6459]<=8'd211;
		data_a[6460]<=8'd211;
		data_a[6461]<=8'd210;
		data_a[6462]<=8'd208;
		data_a[6463]<=8'd208;
		data_a[6464]<=8'd208;
		data_a[6465]<=8'd208;
		data_a[6466]<=8'd206;
		data_a[6467]<=8'd207;
		data_a[6468]<=8'd170;
		data_a[6469]<=8'd189;
		data_a[6470]<=8'd189;
		data_a[6471]<=8'd147;
		data_a[6472]<=8'd150;
		data_a[6473]<=8'd122;
		data_a[6474]<=8'd118;
		data_a[6475]<=8'd127;
		data_a[6476]<=8'd129;
		data_a[6477]<=8'd103;
		data_a[6478]<=8'd81;
		data_a[6479]<=8'd83;
		data_a[6480]<=8'd76;
		data_a[6481]<=8'd77;
		data_a[6482]<=8'd74;
		data_a[6483]<=8'd67;
		data_a[6484]<=8'd77;
		data_a[6485]<=8'd70;
		data_a[6486]<=8'd73;
		data_a[6487]<=8'd69;
		data_a[6488]<=8'd68;
		data_a[6489]<=8'd64;
		data_a[6490]<=8'd61;
		data_a[6491]<=8'd58;
		data_a[6492]<=8'd70;
		data_a[6493]<=8'd59;
		data_a[6494]<=8'd72;
		data_a[6495]<=8'd63;
		data_a[6496]<=8'd72;
		data_a[6497]<=8'd70;
		data_a[6498]<=8'd72;
		data_a[6499]<=8'd77;
		data_a[6500]<=8'd82;
		data_a[6501]<=8'd83;
		data_a[6502]<=8'd81;
		data_a[6503]<=8'd81;
		data_a[6504]<=8'd87;
		data_a[6505]<=8'd91;
		data_a[6506]<=8'd94;
		data_a[6507]<=8'd98;
		data_a[6508]<=8'd91;
		data_a[6509]<=8'd90;
		data_a[6510]<=8'd93;
		data_a[6511]<=8'd87;
		data_a[6512]<=8'd92;
		data_a[6513]<=8'd89;
		data_a[6514]<=8'd91;
		data_a[6515]<=8'd128;
		data_a[6516]<=8'd183;
		data_a[6517]<=8'd203;
		data_a[6518]<=8'd203;
		data_a[6519]<=8'd208;
		data_a[6520]<=8'd212;
		data_a[6521]<=8'd212;
		data_a[6522]<=8'd214;
		data_a[6523]<=8'd205;
		data_a[6524]<=8'd210;
		data_a[6525]<=8'd215;
		data_a[6526]<=8'd195;
		data_a[6527]<=8'd88;
		data_a[6528]<=8'd80;
		data_a[6529]<=8'd73;
		data_a[6530]<=8'd69;
		data_a[6531]<=8'd66;
		data_a[6532]<=8'd66;
		data_a[6533]<=8'd86;
		data_a[6534]<=8'd104;
		data_a[6535]<=8'd117;
		data_a[6536]<=8'd130;
		data_a[6537]<=8'd144;
		data_a[6538]<=8'd145;
		data_a[6539]<=8'd147;
		data_a[6540]<=8'd157;
		data_a[6541]<=8'd160;
		data_a[6542]<=8'd162;
		data_a[6543]<=8'd166;
		data_a[6544]<=8'd164;
		data_a[6545]<=8'd167;
		data_a[6546]<=8'd171;
		data_a[6547]<=8'd171;
		data_a[6548]<=8'd174;
		data_a[6549]<=8'd174;
		data_a[6550]<=8'd171;
		data_a[6551]<=8'd170;
		data_a[6552]<=8'd168;
		data_a[6553]<=8'd163;
		data_a[6554]<=8'd153;
		data_a[6555]<=8'd163;
		data_a[6556]<=8'd173;
		data_a[6557]<=8'd178;
		data_a[6558]<=8'd181;
		data_a[6559]<=8'd182;
		data_a[6560]<=8'd183;
		data_a[6561]<=8'd181;
		data_a[6562]<=8'd179;
		data_a[6563]<=8'd180;
		data_a[6564]<=8'd182;
		data_a[6565]<=8'd181;
		data_a[6566]<=8'd182;
		data_a[6567]<=8'd186;
		data_a[6568]<=8'd184;
		data_a[6569]<=8'd176;
		data_a[6570]<=8'd149;
		data_a[6571]<=8'd119;
		data_a[6572]<=8'd115;
		data_a[6573]<=8'd112;
		data_a[6574]<=8'd128;
		data_a[6575]<=8'd142;
		data_a[6576]<=8'd152;
		data_a[6577]<=8'd215;
		data_a[6578]<=8'd216;
		data_a[6579]<=8'd218;
		data_a[6580]<=8'd219;
		data_a[6581]<=8'd219;
		data_a[6582]<=8'd220;
		data_a[6583]<=8'd222;
		data_a[6584]<=8'd222;
		data_a[6585]<=8'd221;
		data_a[6586]<=8'd223;
		data_a[6587]<=8'd223;
		data_a[6588]<=8'd224;
		data_a[6589]<=8'd226;
		data_a[6590]<=8'd227;
		data_a[6591]<=8'd227;
		data_a[6592]<=8'd228;
		data_a[6593]<=8'd230;
		data_a[6594]<=8'd231;
		data_a[6595]<=8'd232;
		data_a[6596]<=8'd233;
		data_a[6597]<=8'd233;
		data_a[6598]<=8'd233;
		data_a[6599]<=8'd234;
		data_a[6600]<=8'd255;
		data_a[6601]<=8'd217;
		data_a[6602]<=8'd213;
		data_a[6603]<=8'd211;
		data_a[6604]<=8'd207;
		data_a[6605]<=8'd209;
		data_a[6606]<=8'd209;
		data_a[6607]<=8'd213;
		data_a[6608]<=8'd210;
		data_a[6609]<=8'd211;
		data_a[6610]<=8'd211;
		data_a[6611]<=8'd209;
		data_a[6612]<=8'd207;
		data_a[6613]<=8'd207;
		data_a[6614]<=8'd208;
		data_a[6615]<=8'd208;
		data_a[6616]<=8'd202;
		data_a[6617]<=8'd212;
		data_a[6618]<=8'd188;
		data_a[6619]<=8'd191;
		data_a[6620]<=8'd172;
		data_a[6621]<=8'd124;
		data_a[6622]<=8'd97;
		data_a[6623]<=8'd174;
		data_a[6624]<=8'd187;
		data_a[6625]<=8'd173;
		data_a[6626]<=8'd207;
		data_a[6627]<=8'd100;
		data_a[6628]<=8'd83;
		data_a[6629]<=8'd81;
		data_a[6630]<=8'd82;
		data_a[6631]<=8'd77;
		data_a[6632]<=8'd71;
		data_a[6633]<=8'd74;
		data_a[6634]<=8'd71;
		data_a[6635]<=8'd71;
		data_a[6636]<=8'd64;
		data_a[6637]<=8'd68;
		data_a[6638]<=8'd57;
		data_a[6639]<=8'd64;
		data_a[6640]<=8'd61;
		data_a[6641]<=8'd65;
		data_a[6642]<=8'd65;
		data_a[6643]<=8'd74;
		data_a[6644]<=8'd68;
		data_a[6645]<=8'd69;
		data_a[6646]<=8'd70;
		data_a[6647]<=8'd78;
		data_a[6648]<=8'd69;
		data_a[6649]<=8'd73;
		data_a[6650]<=8'd80;
		data_a[6651]<=8'd82;
		data_a[6652]<=8'd80;
		data_a[6653]<=8'd77;
		data_a[6654]<=8'd80;
		data_a[6655]<=8'd88;
		data_a[6656]<=8'd90;
		data_a[6657]<=8'd94;
		data_a[6658]<=8'd89;
		data_a[6659]<=8'd90;
		data_a[6660]<=8'd93;
		data_a[6661]<=8'd100;
		data_a[6662]<=8'd98;
		data_a[6663]<=8'd92;
		data_a[6664]<=8'd105;
		data_a[6665]<=8'd156;
		data_a[6666]<=8'd147;
		data_a[6667]<=8'd205;
		data_a[6668]<=8'd215;
		data_a[6669]<=8'd208;
		data_a[6670]<=8'd205;
		data_a[6671]<=8'd211;
		data_a[6672]<=8'd212;
		data_a[6673]<=8'd212;
		data_a[6674]<=8'd206;
		data_a[6675]<=8'd210;
		data_a[6676]<=8'd196;
		data_a[6677]<=8'd77;
		data_a[6678]<=8'd83;
		data_a[6679]<=8'd71;
		data_a[6680]<=8'd70;
		data_a[6681]<=8'd66;
		data_a[6682]<=8'd72;
		data_a[6683]<=8'd99;
		data_a[6684]<=8'd110;
		data_a[6685]<=8'd126;
		data_a[6686]<=8'd137;
		data_a[6687]<=8'd142;
		data_a[6688]<=8'd147;
		data_a[6689]<=8'd150;
		data_a[6690]<=8'd160;
		data_a[6691]<=8'd162;
		data_a[6692]<=8'd163;
		data_a[6693]<=8'd167;
		data_a[6694]<=8'd165;
		data_a[6695]<=8'd170;
		data_a[6696]<=8'd168;
		data_a[6697]<=8'd168;
		data_a[6698]<=8'd171;
		data_a[6699]<=8'd172;
		data_a[6700]<=8'd172;
		data_a[6701]<=8'd173;
		data_a[6702]<=8'd174;
		data_a[6703]<=8'd171;
		data_a[6704]<=8'd171;
		data_a[6705]<=8'd176;
		data_a[6706]<=8'd180;
		data_a[6707]<=8'd182;
		data_a[6708]<=8'd182;
		data_a[6709]<=8'd184;
		data_a[6710]<=8'd183;
		data_a[6711]<=8'd181;
		data_a[6712]<=8'd180;
		data_a[6713]<=8'd181;
		data_a[6714]<=8'd181;
		data_a[6715]<=8'd181;
		data_a[6716]<=8'd183;
		data_a[6717]<=8'd186;
		data_a[6718]<=8'd184;
		data_a[6719]<=8'd177;
		data_a[6720]<=8'd149;
		data_a[6721]<=8'd119;
		data_a[6722]<=8'd116;
		data_a[6723]<=8'd113;
		data_a[6724]<=8'd123;
		data_a[6725]<=8'd127;
		data_a[6726]<=8'd141;
		data_a[6727]<=8'd210;
		data_a[6728]<=8'd216;
		data_a[6729]<=8'd217;
		data_a[6730]<=8'd217;
		data_a[6731]<=8'd218;
		data_a[6732]<=8'd219;
		data_a[6733]<=8'd221;
		data_a[6734]<=8'd222;
		data_a[6735]<=8'd222;
		data_a[6736]<=8'd222;
		data_a[6737]<=8'd221;
		data_a[6738]<=8'd221;
		data_a[6739]<=8'd223;
		data_a[6740]<=8'd225;
		data_a[6741]<=8'd227;
		data_a[6742]<=8'd230;
		data_a[6743]<=8'd233;
		data_a[6744]<=8'd235;
		data_a[6745]<=8'd235;
		data_a[6746]<=8'd234;
		data_a[6747]<=8'd232;
		data_a[6748]<=8'd232;
		data_a[6749]<=8'd234;
		data_a[6750]<=8'd253;
		data_a[6751]<=8'd202;
		data_a[6752]<=8'd201;
		data_a[6753]<=8'd213;
		data_a[6754]<=8'd210;
		data_a[6755]<=8'd211;
		data_a[6756]<=8'd207;
		data_a[6757]<=8'd208;
		data_a[6758]<=8'd210;
		data_a[6759]<=8'd211;
		data_a[6760]<=8'd210;
		data_a[6761]<=8'd208;
		data_a[6762]<=8'd206;
		data_a[6763]<=8'd207;
		data_a[6764]<=8'd207;
		data_a[6765]<=8'd207;
		data_a[6766]<=8'd209;
		data_a[6767]<=8'd207;
		data_a[6768]<=8'd200;
		data_a[6769]<=8'd151;
		data_a[6770]<=8'd129;
		data_a[6771]<=8'd129;
		data_a[6772]<=8'd182;
		data_a[6773]<=8'd156;
		data_a[6774]<=8'd109;
		data_a[6775]<=8'd99;
		data_a[6776]<=8'd70;
		data_a[6777]<=8'd82;
		data_a[6778]<=8'd84;
		data_a[6779]<=8'd88;
		data_a[6780]<=8'd93;
		data_a[6781]<=8'd80;
		data_a[6782]<=8'd72;
		data_a[6783]<=8'd71;
		data_a[6784]<=8'd69;
		data_a[6785]<=8'd59;
		data_a[6786]<=8'd66;
		data_a[6787]<=8'd60;
		data_a[6788]<=8'd61;
		data_a[6789]<=8'd65;
		data_a[6790]<=8'd60;
		data_a[6791]<=8'd63;
		data_a[6792]<=8'd62;
		data_a[6793]<=8'd73;
		data_a[6794]<=8'd66;
		data_a[6795]<=8'd63;
		data_a[6796]<=8'd65;
		data_a[6797]<=8'd74;
		data_a[6798]<=8'd72;
		data_a[6799]<=8'd72;
		data_a[6800]<=8'd78;
		data_a[6801]<=8'd82;
		data_a[6802]<=8'd83;
		data_a[6803]<=8'd79;
		data_a[6804]<=8'd78;
		data_a[6805]<=8'd88;
		data_a[6806]<=8'd90;
		data_a[6807]<=8'd89;
		data_a[6808]<=8'd91;
		data_a[6809]<=8'd90;
		data_a[6810]<=8'd84;
		data_a[6811]<=8'd101;
		data_a[6812]<=8'd101;
		data_a[6813]<=8'd87;
		data_a[6814]<=8'd102;
		data_a[6815]<=8'd122;
		data_a[6816]<=8'd169;
		data_a[6817]<=8'd182;
		data_a[6818]<=8'd200;
		data_a[6819]<=8'd206;
		data_a[6820]<=8'd216;
		data_a[6821]<=8'd204;
		data_a[6822]<=8'd212;
		data_a[6823]<=8'd207;
		data_a[6824]<=8'd215;
		data_a[6825]<=8'd214;
		data_a[6826]<=8'd178;
		data_a[6827]<=8'd80;
		data_a[6828]<=8'd84;
		data_a[6829]<=8'd74;
		data_a[6830]<=8'd72;
		data_a[6831]<=8'd66;
		data_a[6832]<=8'd81;
		data_a[6833]<=8'd108;
		data_a[6834]<=8'd120;
		data_a[6835]<=8'd137;
		data_a[6836]<=8'd144;
		data_a[6837]<=8'd141;
		data_a[6838]<=8'd151;
		data_a[6839]<=8'd154;
		data_a[6840]<=8'd161;
		data_a[6841]<=8'd163;
		data_a[6842]<=8'd164;
		data_a[6843]<=8'd166;
		data_a[6844]<=8'd167;
		data_a[6845]<=8'd170;
		data_a[6846]<=8'd170;
		data_a[6847]<=8'd170;
		data_a[6848]<=8'd171;
		data_a[6849]<=8'd171;
		data_a[6850]<=8'd171;
		data_a[6851]<=8'd174;
		data_a[6852]<=8'd177;
		data_a[6853]<=8'd177;
		data_a[6854]<=8'd181;
		data_a[6855]<=8'd182;
		data_a[6856]<=8'd181;
		data_a[6857]<=8'd183;
		data_a[6858]<=8'd181;
		data_a[6859]<=8'd184;
		data_a[6860]<=8'd182;
		data_a[6861]<=8'd181;
		data_a[6862]<=8'd182;
		data_a[6863]<=8'd182;
		data_a[6864]<=8'd181;
		data_a[6865]<=8'd180;
		data_a[6866]<=8'd183;
		data_a[6867]<=8'd185;
		data_a[6868]<=8'd182;
		data_a[6869]<=8'd177;
		data_a[6870]<=8'd148;
		data_a[6871]<=8'd134;
		data_a[6872]<=8'd119;
		data_a[6873]<=8'd106;
		data_a[6874]<=8'd123;
		data_a[6875]<=8'd129;
		data_a[6876]<=8'd137;
		data_a[6877]<=8'd216;
		data_a[6878]<=8'd216;
		data_a[6879]<=8'd216;
		data_a[6880]<=8'd216;
		data_a[6881]<=8'd217;
		data_a[6882]<=8'd219;
		data_a[6883]<=8'd220;
		data_a[6884]<=8'd221;
		data_a[6885]<=8'd221;
		data_a[6886]<=8'd221;
		data_a[6887]<=8'd219;
		data_a[6888]<=8'd219;
		data_a[6889]<=8'd223;
		data_a[6890]<=8'd227;
		data_a[6891]<=8'd228;
		data_a[6892]<=8'd229;
		data_a[6893]<=8'd231;
		data_a[6894]<=8'd234;
		data_a[6895]<=8'd236;
		data_a[6896]<=8'd239;
		data_a[6897]<=8'd241;
		data_a[6898]<=8'd243;
		data_a[6899]<=8'd245;
		data_a[6900]<=8'd255;
		data_a[6901]<=8'd188;
		data_a[6902]<=8'd191;
		data_a[6903]<=8'd221;
		data_a[6904]<=8'd215;
		data_a[6905]<=8'd208;
		data_a[6906]<=8'd205;
		data_a[6907]<=8'd208;
		data_a[6908]<=8'd209;
		data_a[6909]<=8'd210;
		data_a[6910]<=8'd209;
		data_a[6911]<=8'd207;
		data_a[6912]<=8'd206;
		data_a[6913]<=8'd207;
		data_a[6914]<=8'd208;
		data_a[6915]<=8'd208;
		data_a[6916]<=8'd206;
		data_a[6917]<=8'd198;
		data_a[6918]<=8'd200;
		data_a[6919]<=8'd173;
		data_a[6920]<=8'd130;
		data_a[6921]<=8'd142;
		data_a[6922]<=8'd102;
		data_a[6923]<=8'd96;
		data_a[6924]<=8'd73;
		data_a[6925]<=8'd98;
		data_a[6926]<=8'd87;
		data_a[6927]<=8'd86;
		data_a[6928]<=8'd80;
		data_a[6929]<=8'd94;
		data_a[6930]<=8'd181;
		data_a[6931]<=8'd168;
		data_a[6932]<=8'd72;
		data_a[6933]<=8'd70;
		data_a[6934]<=8'd62;
		data_a[6935]<=8'd65;
		data_a[6936]<=8'd64;
		data_a[6937]<=8'd65;
		data_a[6938]<=8'd60;
		data_a[6939]<=8'd59;
		data_a[6940]<=8'd61;
		data_a[6941]<=8'd68;
		data_a[6942]<=8'd58;
		data_a[6943]<=8'd77;
		data_a[6944]<=8'd61;
		data_a[6945]<=8'd67;
		data_a[6946]<=8'd62;
		data_a[6947]<=8'd71;
		data_a[6948]<=8'd69;
		data_a[6949]<=8'd68;
		data_a[6950]<=8'd72;
		data_a[6951]<=8'd77;
		data_a[6952]<=8'd82;
		data_a[6953]<=8'd82;
		data_a[6954]<=8'd81;
		data_a[6955]<=8'd91;
		data_a[6956]<=8'd88;
		data_a[6957]<=8'd87;
		data_a[6958]<=8'd88;
		data_a[6959]<=8'd87;
		data_a[6960]<=8'd83;
		data_a[6961]<=8'd94;
		data_a[6962]<=8'd101;
		data_a[6963]<=8'd94;
		data_a[6964]<=8'd93;
		data_a[6965]<=8'd118;
		data_a[6966]<=8'd135;
		data_a[6967]<=8'd168;
		data_a[6968]<=8'd207;
		data_a[6969]<=8'd209;
		data_a[6970]<=8'd205;
		data_a[6971]<=8'd210;
		data_a[6972]<=8'd207;
		data_a[6973]<=8'd212;
		data_a[6974]<=8'd210;
		data_a[6975]<=8'd203;
		data_a[6976]<=8'd195;
		data_a[6977]<=8'd78;
		data_a[6978]<=8'd84;
		data_a[6979]<=8'd68;
		data_a[6980]<=8'd70;
		data_a[6981]<=8'd67;
		data_a[6982]<=8'd94;
		data_a[6983]<=8'd117;
		data_a[6984]<=8'd136;
		data_a[6985]<=8'd143;
		data_a[6986]<=8'd147;
		data_a[6987]<=8'd146;
		data_a[6988]<=8'd153;
		data_a[6989]<=8'd157;
		data_a[6990]<=8'd159;
		data_a[6991]<=8'd163;
		data_a[6992]<=8'd165;
		data_a[6993]<=8'd165;
		data_a[6994]<=8'd168;
		data_a[6995]<=8'd169;
		data_a[6996]<=8'd171;
		data_a[6997]<=8'd170;
		data_a[6998]<=8'd171;
		data_a[6999]<=8'd170;
		data_a[7000]<=8'd168;
		data_a[7001]<=8'd170;
		data_a[7002]<=8'd174;
		data_a[7003]<=8'd174;
		data_a[7004]<=8'd180;
		data_a[7005]<=8'd181;
		data_a[7006]<=8'd178;
		data_a[7007]<=8'd182;
		data_a[7008]<=8'd179;
		data_a[7009]<=8'd182;
		data_a[7010]<=8'd180;
		data_a[7011]<=8'd183;
		data_a[7012]<=8'd184;
		data_a[7013]<=8'd185;
		data_a[7014]<=8'd184;
		data_a[7015]<=8'd184;
		data_a[7016]<=8'd186;
		data_a[7017]<=8'd186;
		data_a[7018]<=8'd181;
		data_a[7019]<=8'd177;
		data_a[7020]<=8'd163;
		data_a[7021]<=8'd124;
		data_a[7022]<=8'd116;
		data_a[7023]<=8'd116;
		data_a[7024]<=8'd119;
		data_a[7025]<=8'd129;
		data_a[7026]<=8'd139;
		data_a[7027]<=8'd217;
		data_a[7028]<=8'd216;
		data_a[7029]<=8'd215;
		data_a[7030]<=8'd215;
		data_a[7031]<=8'd218;
		data_a[7032]<=8'd220;
		data_a[7033]<=8'd220;
		data_a[7034]<=8'd219;
		data_a[7035]<=8'd219;
		data_a[7036]<=8'd219;
		data_a[7037]<=8'd219;
		data_a[7038]<=8'd220;
		data_a[7039]<=8'd224;
		data_a[7040]<=8'd227;
		data_a[7041]<=8'd229;
		data_a[7042]<=8'd233;
		data_a[7043]<=8'd238;
		data_a[7044]<=8'd242;
		data_a[7045]<=8'd246;
		data_a[7046]<=8'd250;
		data_a[7047]<=8'd253;
		data_a[7048]<=8'd255;
		data_a[7049]<=8'd255;
		data_a[7050]<=8'd254;
		data_a[7051]<=8'd214;
		data_a[7052]<=8'd211;
		data_a[7053]<=8'd211;
		data_a[7054]<=8'd203;
		data_a[7055]<=8'd213;
		data_a[7056]<=8'd211;
		data_a[7057]<=8'd208;
		data_a[7058]<=8'd207;
		data_a[7059]<=8'd208;
		data_a[7060]<=8'd208;
		data_a[7061]<=8'd206;
		data_a[7062]<=8'd206;
		data_a[7063]<=8'd208;
		data_a[7064]<=8'd210;
		data_a[7065]<=8'd210;
		data_a[7066]<=8'd196;
		data_a[7067]<=8'd192;
		data_a[7068]<=8'd190;
		data_a[7069]<=8'd164;
		data_a[7070]<=8'd115;
		data_a[7071]<=8'd85;
		data_a[7072]<=8'd115;
		data_a[7073]<=8'd113;
		data_a[7074]<=8'd202;
		data_a[7075]<=8'd179;
		data_a[7076]<=8'd115;
		data_a[7077]<=8'd146;
		data_a[7078]<=8'd208;
		data_a[7079]<=8'd156;
		data_a[7080]<=8'd213;
		data_a[7081]<=8'd123;
		data_a[7082]<=8'd88;
		data_a[7083]<=8'd75;
		data_a[7084]<=8'd62;
		data_a[7085]<=8'd61;
		data_a[7086]<=8'd60;
		data_a[7087]<=8'd59;
		data_a[7088]<=8'd63;
		data_a[7089]<=8'd54;
		data_a[7090]<=8'd60;
		data_a[7091]<=8'd62;
		data_a[7092]<=8'd59;
		data_a[7093]<=8'd65;
		data_a[7094]<=8'd63;
		data_a[7095]<=8'd60;
		data_a[7096]<=8'd62;
		data_a[7097]<=8'd63;
		data_a[7098]<=8'd71;
		data_a[7099]<=8'd67;
		data_a[7100]<=8'd68;
		data_a[7101]<=8'd69;
		data_a[7102]<=8'd76;
		data_a[7103]<=8'd77;
		data_a[7104]<=8'd74;
		data_a[7105]<=8'd82;
		data_a[7106]<=8'd86;
		data_a[7107]<=8'd84;
		data_a[7108]<=8'd78;
		data_a[7109]<=8'd80;
		data_a[7110]<=8'd90;
		data_a[7111]<=8'd84;
		data_a[7112]<=8'd89;
		data_a[7113]<=8'd92;
		data_a[7114]<=8'd106;
		data_a[7115]<=8'd109;
		data_a[7116]<=8'd130;
		data_a[7117]<=8'd153;
		data_a[7118]<=8'd202;
		data_a[7119]<=8'd205;
		data_a[7120]<=8'd198;
		data_a[7121]<=8'd204;
		data_a[7122]<=8'd200;
		data_a[7123]<=8'd212;
		data_a[7124]<=8'd207;
		data_a[7125]<=8'd217;
		data_a[7126]<=8'd189;
		data_a[7127]<=8'd83;
		data_a[7128]<=8'd71;
		data_a[7129]<=8'd71;
		data_a[7130]<=8'd64;
		data_a[7131]<=8'd67;
		data_a[7132]<=8'd106;
		data_a[7133]<=8'd124;
		data_a[7134]<=8'd149;
		data_a[7135]<=8'd145;
		data_a[7136]<=8'd147;
		data_a[7137]<=8'd152;
		data_a[7138]<=8'd155;
		data_a[7139]<=8'd158;
		data_a[7140]<=8'd157;
		data_a[7141]<=8'd162;
		data_a[7142]<=8'd165;
		data_a[7143]<=8'd165;
		data_a[7144]<=8'd170;
		data_a[7145]<=8'd169;
		data_a[7146]<=8'd169;
		data_a[7147]<=8'd170;
		data_a[7148]<=8'd172;
		data_a[7149]<=8'd173;
		data_a[7150]<=8'd172;
		data_a[7151]<=8'd174;
		data_a[7152]<=8'd177;
		data_a[7153]<=8'd177;
		data_a[7154]<=8'd178;
		data_a[7155]<=8'd179;
		data_a[7156]<=8'd178;
		data_a[7157]<=8'd182;
		data_a[7158]<=8'd178;
		data_a[7159]<=8'd180;
		data_a[7160]<=8'd179;
		data_a[7161]<=8'd183;
		data_a[7162]<=8'd185;
		data_a[7163]<=8'd188;
		data_a[7164]<=8'd189;
		data_a[7165]<=8'd189;
		data_a[7166]<=8'd191;
		data_a[7167]<=8'd188;
		data_a[7168]<=8'd181;
		data_a[7169]<=8'd177;
		data_a[7170]<=8'd158;
		data_a[7171]<=8'd125;
		data_a[7172]<=8'd117;
		data_a[7173]<=8'd111;
		data_a[7174]<=8'd116;
		data_a[7175]<=8'd117;
		data_a[7176]<=8'd141;
		data_a[7177]<=8'd203;
		data_a[7178]<=8'd215;
		data_a[7179]<=8'd214;
		data_a[7180]<=8'd215;
		data_a[7181]<=8'd219;
		data_a[7182]<=8'd220;
		data_a[7183]<=8'd219;
		data_a[7184]<=8'd218;
		data_a[7185]<=8'd217;
		data_a[7186]<=8'd220;
		data_a[7187]<=8'd220;
		data_a[7188]<=8'd222;
		data_a[7189]<=8'd222;
		data_a[7190]<=8'd222;
		data_a[7191]<=8'd228;
		data_a[7192]<=8'd242;
		data_a[7193]<=8'd255;
		data_a[7194]<=8'd253;
		data_a[7195]<=8'd253;
		data_a[7196]<=8'd253;
		data_a[7197]<=8'd252;
		data_a[7198]<=8'd253;
		data_a[7199]<=8'd254;
		data_a[7200]<=8'd254;
		data_a[7201]<=8'd213;
		data_a[7202]<=8'd216;
		data_a[7203]<=8'd216;
		data_a[7204]<=8'd204;
		data_a[7205]<=8'd202;
		data_a[7206]<=8'd204;
		data_a[7207]<=8'd208;
		data_a[7208]<=8'd206;
		data_a[7209]<=8'd212;
		data_a[7210]<=8'd207;
		data_a[7211]<=8'd207;
		data_a[7212]<=8'd215;
		data_a[7213]<=8'd207;
		data_a[7214]<=8'd172;
		data_a[7215]<=8'd200;
		data_a[7216]<=8'd207;
		data_a[7217]<=8'd204;
		data_a[7218]<=8'd191;
		data_a[7219]<=8'd115;
		data_a[7220]<=8'd158;
		data_a[7221]<=8'd217;
		data_a[7222]<=8'd125;
		data_a[7223]<=8'd122;
		data_a[7224]<=8'd121;
		data_a[7225]<=8'd125;
		data_a[7226]<=8'd76;
		data_a[7227]<=8'd201;
		data_a[7228]<=8'd250;
		data_a[7229]<=8'd185;
		data_a[7230]<=8'd222;
		data_a[7231]<=8'd120;
		data_a[7232]<=8'd94;
		data_a[7233]<=8'd71;
		data_a[7234]<=8'd60;
		data_a[7235]<=8'd58;
		data_a[7236]<=8'd61;
		data_a[7237]<=8'd64;
		data_a[7238]<=8'd60;
		data_a[7239]<=8'd59;
		data_a[7240]<=8'd62;
		data_a[7241]<=8'd61;
		data_a[7242]<=8'd62;
		data_a[7243]<=8'd63;
		data_a[7244]<=8'd65;
		data_a[7245]<=8'd65;
		data_a[7246]<=8'd63;
		data_a[7247]<=8'd61;
		data_a[7248]<=8'd70;
		data_a[7249]<=8'd72;
		data_a[7250]<=8'd69;
		data_a[7251]<=8'd66;
		data_a[7252]<=8'd79;
		data_a[7253]<=8'd74;
		data_a[7254]<=8'd72;
		data_a[7255]<=8'd76;
		data_a[7256]<=8'd79;
		data_a[7257]<=8'd75;
		data_a[7258]<=8'd76;
		data_a[7259]<=8'd77;
		data_a[7260]<=8'd86;
		data_a[7261]<=8'd84;
		data_a[7262]<=8'd84;
		data_a[7263]<=8'd85;
		data_a[7264]<=8'd102;
		data_a[7265]<=8'd115;
		data_a[7266]<=8'd141;
		data_a[7267]<=8'd162;
		data_a[7268]<=8'd175;
		data_a[7269]<=8'd175;
		data_a[7270]<=8'd194;
		data_a[7271]<=8'd201;
		data_a[7272]<=8'd212;
		data_a[7273]<=8'd206;
		data_a[7274]<=8'd212;
		data_a[7275]<=8'd215;
		data_a[7276]<=8'd185;
		data_a[7277]<=8'd84;
		data_a[7278]<=8'd77;
		data_a[7279]<=8'd68;
		data_a[7280]<=8'd69;
		data_a[7281]<=8'd81;
		data_a[7282]<=8'd113;
		data_a[7283]<=8'd126;
		data_a[7284]<=8'd146;
		data_a[7285]<=8'd150;
		data_a[7286]<=8'd153;
		data_a[7287]<=8'd153;
		data_a[7288]<=8'd157;
		data_a[7289]<=8'd158;
		data_a[7290]<=8'd162;
		data_a[7291]<=8'd166;
		data_a[7292]<=8'd167;
		data_a[7293]<=8'd166;
		data_a[7294]<=8'd168;
		data_a[7295]<=8'd171;
		data_a[7296]<=8'd170;
		data_a[7297]<=8'd170;
		data_a[7298]<=8'd175;
		data_a[7299]<=8'd177;
		data_a[7300]<=8'd173;
		data_a[7301]<=8'd179;
		data_a[7302]<=8'd173;
		data_a[7303]<=8'd175;
		data_a[7304]<=8'd183;
		data_a[7305]<=8'd175;
		data_a[7306]<=8'd176;
		data_a[7307]<=8'd177;
		data_a[7308]<=8'd174;
		data_a[7309]<=8'd178;
		data_a[7310]<=8'd178;
		data_a[7311]<=8'd185;
		data_a[7312]<=8'd184;
		data_a[7313]<=8'd191;
		data_a[7314]<=8'd191;
		data_a[7315]<=8'd195;
		data_a[7316]<=8'd192;
		data_a[7317]<=8'd187;
		data_a[7318]<=8'd185;
		data_a[7319]<=8'd182;
		data_a[7320]<=8'd168;
		data_a[7321]<=8'd144;
		data_a[7322]<=8'd116;
		data_a[7323]<=8'd111;
		data_a[7324]<=8'd122;
		data_a[7325]<=8'd126;
		data_a[7326]<=8'd138;
		data_a[7327]<=8'd193;
		data_a[7328]<=8'd214;
		data_a[7329]<=8'd215;
		data_a[7330]<=8'd216;
		data_a[7331]<=8'd218;
		data_a[7332]<=8'd219;
		data_a[7333]<=8'd219;
		data_a[7334]<=8'd218;
		data_a[7335]<=8'd217;
		data_a[7336]<=8'd221;
		data_a[7337]<=8'd222;
		data_a[7338]<=8'd218;
		data_a[7339]<=8'd220;
		data_a[7340]<=8'd246;
		data_a[7341]<=8'd252;
		data_a[7342]<=8'd254;
		data_a[7343]<=8'd255;
		data_a[7344]<=8'd255;
		data_a[7345]<=8'd255;
		data_a[7346]<=8'd255;
		data_a[7347]<=8'd255;
		data_a[7348]<=8'd255;
		data_a[7349]<=8'd255;
		data_a[7350]<=8'd255;
		data_a[7351]<=8'd212;
		data_a[7352]<=8'd210;
		data_a[7353]<=8'd215;
		data_a[7354]<=8'd219;
		data_a[7355]<=8'd216;
		data_a[7356]<=8'd204;
		data_a[7357]<=8'd199;
		data_a[7358]<=8'd212;
		data_a[7359]<=8'd211;
		data_a[7360]<=8'd207;
		data_a[7361]<=8'd190;
		data_a[7362]<=8'd198;
		data_a[7363]<=8'd198;
		data_a[7364]<=8'd201;
		data_a[7365]<=8'd211;
		data_a[7366]<=8'd204;
		data_a[7367]<=8'd208;
		data_a[7368]<=8'd179;
		data_a[7369]<=8'd192;
		data_a[7370]<=8'd169;
		data_a[7371]<=8'd152;
		data_a[7372]<=8'd150;
		data_a[7373]<=8'd128;
		data_a[7374]<=8'd117;
		data_a[7375]<=8'd104;
		data_a[7376]<=8'd153;
		data_a[7377]<=8'd149;
		data_a[7378]<=8'd114;
		data_a[7379]<=8'd118;
		data_a[7380]<=8'd88;
		data_a[7381]<=8'd68;
		data_a[7382]<=8'd69;
		data_a[7383]<=8'd64;
		data_a[7384]<=8'd58;
		data_a[7385]<=8'd62;
		data_a[7386]<=8'd66;
		data_a[7387]<=8'd61;
		data_a[7388]<=8'd60;
		data_a[7389]<=8'd63;
		data_a[7390]<=8'd62;
		data_a[7391]<=8'd60;
		data_a[7392]<=8'd61;
		data_a[7393]<=8'd65;
		data_a[7394]<=8'd65;
		data_a[7395]<=8'd62;
		data_a[7396]<=8'd63;
		data_a[7397]<=8'd68;
		data_a[7398]<=8'd68;
		data_a[7399]<=8'd68;
		data_a[7400]<=8'd70;
		data_a[7401]<=8'd69;
		data_a[7402]<=8'd76;
		data_a[7403]<=8'd72;
		data_a[7404]<=8'd73;
		data_a[7405]<=8'd74;
		data_a[7406]<=8'd75;
		data_a[7407]<=8'd75;
		data_a[7408]<=8'd74;
		data_a[7409]<=8'd77;
		data_a[7410]<=8'd80;
		data_a[7411]<=8'd81;
		data_a[7412]<=8'd81;
		data_a[7413]<=8'd85;
		data_a[7414]<=8'd94;
		data_a[7415]<=8'd118;
		data_a[7416]<=8'd150;
		data_a[7417]<=8'd122;
		data_a[7418]<=8'd170;
		data_a[7419]<=8'd182;
		data_a[7420]<=8'd175;
		data_a[7421]<=8'd194;
		data_a[7422]<=8'd204;
		data_a[7423]<=8'd208;
		data_a[7424]<=8'd205;
		data_a[7425]<=8'd207;
		data_a[7426]<=8'd199;
		data_a[7427]<=8'd86;
		data_a[7428]<=8'd70;
		data_a[7429]<=8'd64;
		data_a[7430]<=8'd65;
		data_a[7431]<=8'd87;
		data_a[7432]<=8'd121;
		data_a[7433]<=8'd132;
		data_a[7434]<=8'd146;
		data_a[7435]<=8'd146;
		data_a[7436]<=8'd149;
		data_a[7437]<=8'd153;
		data_a[7438]<=8'd157;
		data_a[7439]<=8'd161;
		data_a[7440]<=8'd164;
		data_a[7441]<=8'd166;
		data_a[7442]<=8'd167;
		data_a[7443]<=8'd169;
		data_a[7444]<=8'd171;
		data_a[7445]<=8'd172;
		data_a[7446]<=8'd170;
		data_a[7447]<=8'd174;
		data_a[7448]<=8'd176;
		data_a[7449]<=8'd176;
		data_a[7450]<=8'd177;
		data_a[7451]<=8'd178;
		data_a[7452]<=8'd179;
		data_a[7453]<=8'd177;
		data_a[7454]<=8'd180;
		data_a[7455]<=8'd174;
		data_a[7456]<=8'd171;
		data_a[7457]<=8'd170;
		data_a[7458]<=8'd177;
		data_a[7459]<=8'd175;
		data_a[7460]<=8'd176;
		data_a[7461]<=8'd179;
		data_a[7462]<=8'd181;
		data_a[7463]<=8'd189;
		data_a[7464]<=8'd190;
		data_a[7465]<=8'd193;
		data_a[7466]<=8'd195;
		data_a[7467]<=8'd201;
		data_a[7468]<=8'd188;
		data_a[7469]<=8'd187;
		data_a[7470]<=8'd170;
		data_a[7471]<=8'd149;
		data_a[7472]<=8'd115;
		data_a[7473]<=8'd112;
		data_a[7474]<=8'd118;
		data_a[7475]<=8'd123;
		data_a[7476]<=8'd139;
		data_a[7477]<=8'd185;
		data_a[7478]<=8'd212;
		data_a[7479]<=8'd215;
		data_a[7480]<=8'd216;
		data_a[7481]<=8'd216;
		data_a[7482]<=8'd216;
		data_a[7483]<=8'd217;
		data_a[7484]<=8'd216;
		data_a[7485]<=8'd214;
		data_a[7486]<=8'd218;
		data_a[7487]<=8'd217;
		data_a[7488]<=8'd221;
		data_a[7489]<=8'd221;
		data_a[7490]<=8'd251;
		data_a[7491]<=8'd255;
		data_a[7492]<=8'd255;
		data_a[7493]<=8'd252;
		data_a[7494]<=8'd254;
		data_a[7495]<=8'd254;
		data_a[7496]<=8'd255;
		data_a[7497]<=8'd255;
		data_a[7498]<=8'd255;
		data_a[7499]<=8'd255;
		data_a[7500]<=8'd254;
		data_a[7501]<=8'd218;
		data_a[7502]<=8'd215;
		data_a[7503]<=8'd213;
		data_a[7504]<=8'd213;
		data_a[7505]<=8'd211;
		data_a[7506]<=8'd207;
		data_a[7507]<=8'd215;
		data_a[7508]<=8'd186;
		data_a[7509]<=8'd192;
		data_a[7510]<=8'd205;
		data_a[7511]<=8'd212;
		data_a[7512]<=8'd216;
		data_a[7513]<=8'd202;
		data_a[7514]<=8'd210;
		data_a[7515]<=8'd202;
		data_a[7516]<=8'd201;
		data_a[7517]<=8'd201;
		data_a[7518]<=8'd190;
		data_a[7519]<=8'd182;
		data_a[7520]<=8'd194;
		data_a[7521]<=8'd117;
		data_a[7522]<=8'd168;
		data_a[7523]<=8'd184;
		data_a[7524]<=8'd151;
		data_a[7525]<=8'd101;
		data_a[7526]<=8'd101;
		data_a[7527]<=8'd116;
		data_a[7528]<=8'd249;
		data_a[7529]<=8'd126;
		data_a[7530]<=8'd74;
		data_a[7531]<=8'd108;
		data_a[7532]<=8'd99;
		data_a[7533]<=8'd67;
		data_a[7534]<=8'd56;
		data_a[7535]<=8'd50;
		data_a[7536]<=8'd52;
		data_a[7537]<=8'd63;
		data_a[7538]<=8'd60;
		data_a[7539]<=8'd58;
		data_a[7540]<=8'd57;
		data_a[7541]<=8'd55;
		data_a[7542]<=8'd57;
		data_a[7543]<=8'd62;
		data_a[7544]<=8'd63;
		data_a[7545]<=8'd61;
		data_a[7546]<=8'd61;
		data_a[7547]<=8'd65;
		data_a[7548]<=8'd66;
		data_a[7549]<=8'd64;
		data_a[7550]<=8'd69;
		data_a[7551]<=8'd72;
		data_a[7552]<=8'd72;
		data_a[7553]<=8'd71;
		data_a[7554]<=8'd74;
		data_a[7555]<=8'd71;
		data_a[7556]<=8'd70;
		data_a[7557]<=8'd73;
		data_a[7558]<=8'd71;
		data_a[7559]<=8'd74;
		data_a[7560]<=8'd72;
		data_a[7561]<=8'd74;
		data_a[7562]<=8'd73;
		data_a[7563]<=8'd79;
		data_a[7564]<=8'd94;
		data_a[7565]<=8'd109;
		data_a[7566]<=8'd122;
		data_a[7567]<=8'd108;
		data_a[7568]<=8'd164;
		data_a[7569]<=8'd170;
		data_a[7570]<=8'd146;
		data_a[7571]<=8'd207;
		data_a[7572]<=8'd206;
		data_a[7573]<=8'd203;
		data_a[7574]<=8'd209;
		data_a[7575]<=8'd209;
		data_a[7576]<=8'd198;
		data_a[7577]<=8'd84;
		data_a[7578]<=8'd69;
		data_a[7579]<=8'd62;
		data_a[7580]<=8'd66;
		data_a[7581]<=8'd95;
		data_a[7582]<=8'd125;
		data_a[7583]<=8'd131;
		data_a[7584]<=8'd143;
		data_a[7585]<=8'd145;
		data_a[7586]<=8'd152;
		data_a[7587]<=8'd160;
		data_a[7588]<=8'd160;
		data_a[7589]<=8'd164;
		data_a[7590]<=8'd167;
		data_a[7591]<=8'd167;
		data_a[7592]<=8'd168;
		data_a[7593]<=8'd172;
		data_a[7594]<=8'd174;
		data_a[7595]<=8'd174;
		data_a[7596]<=8'd170;
		data_a[7597]<=8'd177;
		data_a[7598]<=8'd174;
		data_a[7599]<=8'd172;
		data_a[7600]<=8'd179;
		data_a[7601]<=8'd174;
		data_a[7602]<=8'd178;
		data_a[7603]<=8'd172;
		data_a[7604]<=8'd171;
		data_a[7605]<=8'd170;
		data_a[7606]<=8'd167;
		data_a[7607]<=8'd158;
		data_a[7608]<=8'd167;
		data_a[7609]<=8'd158;
		data_a[7610]<=8'd162;
		data_a[7611]<=8'd165;
		data_a[7612]<=8'd177;
		data_a[7613]<=8'd164;
		data_a[7614]<=8'd175;
		data_a[7615]<=8'd200;
		data_a[7616]<=8'd193;
		data_a[7617]<=8'd189;
		data_a[7618]<=8'd191;
		data_a[7619]<=8'd185;
		data_a[7620]<=8'd175;
		data_a[7621]<=8'd159;
		data_a[7622]<=8'd120;
		data_a[7623]<=8'd113;
		data_a[7624]<=8'd115;
		data_a[7625]<=8'd120;
		data_a[7626]<=8'd138;
		data_a[7627]<=8'd174;
		data_a[7628]<=8'd211;
		data_a[7629]<=8'd215;
		data_a[7630]<=8'd216;
		data_a[7631]<=8'd215;
		data_a[7632]<=8'd214;
		data_a[7633]<=8'd216;
		data_a[7634]<=8'd217;
		data_a[7635]<=8'd215;
		data_a[7636]<=8'd216;
		data_a[7637]<=8'd221;
		data_a[7638]<=8'd219;
		data_a[7639]<=8'd228;
		data_a[7640]<=8'd233;
		data_a[7641]<=8'd255;
		data_a[7642]<=8'd253;
		data_a[7643]<=8'd254;
		data_a[7644]<=8'd255;
		data_a[7645]<=8'd255;
		data_a[7646]<=8'd255;
		data_a[7647]<=8'd255;
		data_a[7648]<=8'd254;
		data_a[7649]<=8'd254;
		data_a[7650]<=8'd253;
		data_a[7651]<=8'd217;
		data_a[7652]<=8'd216;
		data_a[7653]<=8'd215;
		data_a[7654]<=8'd213;
		data_a[7655]<=8'd212;
		data_a[7656]<=8'd210;
		data_a[7657]<=8'd215;
		data_a[7658]<=8'd217;
		data_a[7659]<=8'd195;
		data_a[7660]<=8'd207;
		data_a[7661]<=8'd202;
		data_a[7662]<=8'd212;
		data_a[7663]<=8'd207;
		data_a[7664]<=8'd203;
		data_a[7665]<=8'd203;
		data_a[7666]<=8'd196;
		data_a[7667]<=8'd205;
		data_a[7668]<=8'd194;
		data_a[7669]<=8'd176;
		data_a[7670]<=8'd195;
		data_a[7671]<=8'd143;
		data_a[7672]<=8'd189;
		data_a[7673]<=8'd204;
		data_a[7674]<=8'd141;
		data_a[7675]<=8'd96;
		data_a[7676]<=8'd99;
		data_a[7677]<=8'd119;
		data_a[7678]<=8'd104;
		data_a[7679]<=8'd80;
		data_a[7680]<=8'd66;
		data_a[7681]<=8'd65;
		data_a[7682]<=8'd65;
		data_a[7683]<=8'd66;
		data_a[7684]<=8'd58;
		data_a[7685]<=8'd61;
		data_a[7686]<=8'd64;
		data_a[7687]<=8'd57;
		data_a[7688]<=8'd58;
		data_a[7689]<=8'd61;
		data_a[7690]<=8'd62;
		data_a[7691]<=8'd63;
		data_a[7692]<=8'd62;
		data_a[7693]<=8'd63;
		data_a[7694]<=8'd66;
		data_a[7695]<=8'd69;
		data_a[7696]<=8'd68;
		data_a[7697]<=8'd65;
		data_a[7698]<=8'd63;
		data_a[7699]<=8'd62;
		data_a[7700]<=8'd67;
		data_a[7701]<=8'd70;
		data_a[7702]<=8'd70;
		data_a[7703]<=8'd70;
		data_a[7704]<=8'd71;
		data_a[7705]<=8'd68;
		data_a[7706]<=8'd73;
		data_a[7707]<=8'd75;
		data_a[7708]<=8'd72;
		data_a[7709]<=8'd73;
		data_a[7710]<=8'd72;
		data_a[7711]<=8'd72;
		data_a[7712]<=8'd72;
		data_a[7713]<=8'd77;
		data_a[7714]<=8'd85;
		data_a[7715]<=8'd94;
		data_a[7716]<=8'd108;
		data_a[7717]<=8'd111;
		data_a[7718]<=8'd117;
		data_a[7719]<=8'd113;
		data_a[7720]<=8'd138;
		data_a[7721]<=8'd150;
		data_a[7722]<=8'd203;
		data_a[7723]<=8'd205;
		data_a[7724]<=8'd209;
		data_a[7725]<=8'd205;
		data_a[7726]<=8'd215;
		data_a[7727]<=8'd99;
		data_a[7728]<=8'd61;
		data_a[7729]<=8'd66;
		data_a[7730]<=8'd62;
		data_a[7731]<=8'd98;
		data_a[7732]<=8'd129;
		data_a[7733]<=8'd137;
		data_a[7734]<=8'd151;
		data_a[7735]<=8'd152;
		data_a[7736]<=8'd154;
		data_a[7737]<=8'd159;
		data_a[7738]<=8'd164;
		data_a[7739]<=8'd166;
		data_a[7740]<=8'd167;
		data_a[7741]<=8'd167;
		data_a[7742]<=8'd168;
		data_a[7743]<=8'd171;
		data_a[7744]<=8'd174;
		data_a[7745]<=8'd175;
		data_a[7746]<=8'd174;
		data_a[7747]<=8'd180;
		data_a[7748]<=8'd175;
		data_a[7749]<=8'd173;
		data_a[7750]<=8'd179;
		data_a[7751]<=8'd172;
		data_a[7752]<=8'd169;
		data_a[7753]<=8'd166;
		data_a[7754]<=8'd167;
		data_a[7755]<=8'd158;
		data_a[7756]<=8'd151;
		data_a[7757]<=8'd139;
		data_a[7758]<=8'd141;
		data_a[7759]<=8'd135;
		data_a[7760]<=8'd133;
		data_a[7761]<=8'd131;
		data_a[7762]<=8'd119;
		data_a[7763]<=8'd133;
		data_a[7764]<=8'd135;
		data_a[7765]<=8'd150;
		data_a[7766]<=8'd188;
		data_a[7767]<=8'd201;
		data_a[7768]<=8'd195;
		data_a[7769]<=8'd190;
		data_a[7770]<=8'd181;
		data_a[7771]<=8'd169;
		data_a[7772]<=8'd133;
		data_a[7773]<=8'd113;
		data_a[7774]<=8'd115;
		data_a[7775]<=8'd118;
		data_a[7776]<=8'd132;
		data_a[7777]<=8'd163;
		data_a[7778]<=8'd212;
		data_a[7779]<=8'd213;
		data_a[7780]<=8'd214;
		data_a[7781]<=8'd214;
		data_a[7782]<=8'd215;
		data_a[7783]<=8'd216;
		data_a[7784]<=8'd217;
		data_a[7785]<=8'd217;
		data_a[7786]<=8'd219;
		data_a[7787]<=8'd220;
		data_a[7788]<=8'd223;
		data_a[7789]<=8'd223;
		data_a[7790]<=8'd226;
		data_a[7791]<=8'd252;
		data_a[7792]<=8'd255;
		data_a[7793]<=8'd255;
		data_a[7794]<=8'd254;
		data_a[7795]<=8'd254;
		data_a[7796]<=8'd255;
		data_a[7797]<=8'd255;
		data_a[7798]<=8'd255;
		data_a[7799]<=8'd255;
		data_a[7800]<=8'd255;
		data_a[7801]<=8'd212;
		data_a[7802]<=8'd213;
		data_a[7803]<=8'd216;
		data_a[7804]<=8'd214;
		data_a[7805]<=8'd216;
		data_a[7806]<=8'd212;
		data_a[7807]<=8'd209;
		data_a[7808]<=8'd214;
		data_a[7809]<=8'd208;
		data_a[7810]<=8'd209;
		data_a[7811]<=8'd194;
		data_a[7812]<=8'd203;
		data_a[7813]<=8'd200;
		data_a[7814]<=8'd208;
		data_a[7815]<=8'd205;
		data_a[7816]<=8'd202;
		data_a[7817]<=8'd203;
		data_a[7818]<=8'd208;
		data_a[7819]<=8'd174;
		data_a[7820]<=8'd194;
		data_a[7821]<=8'd155;
		data_a[7822]<=8'd178;
		data_a[7823]<=8'd173;
		data_a[7824]<=8'd140;
		data_a[7825]<=8'd93;
		data_a[7826]<=8'd87;
		data_a[7827]<=8'd92;
		data_a[7828]<=8'd69;
		data_a[7829]<=8'd68;
		data_a[7830]<=8'd77;
		data_a[7831]<=8'd64;
		data_a[7832]<=8'd77;
		data_a[7833]<=8'd55;
		data_a[7834]<=8'd60;
		data_a[7835]<=8'd60;
		data_a[7836]<=8'd58;
		data_a[7837]<=8'd66;
		data_a[7838]<=8'd62;
		data_a[7839]<=8'd61;
		data_a[7840]<=8'd64;
		data_a[7841]<=8'd66;
		data_a[7842]<=8'd66;
		data_a[7843]<=8'd65;
		data_a[7844]<=8'd66;
		data_a[7845]<=8'd69;
		data_a[7846]<=8'd70;
		data_a[7847]<=8'd68;
		data_a[7848]<=8'd67;
		data_a[7849]<=8'd70;
		data_a[7850]<=8'd69;
		data_a[7851]<=8'd71;
		data_a[7852]<=8'd75;
		data_a[7853]<=8'd75;
		data_a[7854]<=8'd71;
		data_a[7855]<=8'd71;
		data_a[7856]<=8'd72;
		data_a[7857]<=8'd71;
		data_a[7858]<=8'd71;
		data_a[7859]<=8'd69;
		data_a[7860]<=8'd73;
		data_a[7861]<=8'd71;
		data_a[7862]<=8'd73;
		data_a[7863]<=8'd74;
		data_a[7864]<=8'd75;
		data_a[7865]<=8'd91;
		data_a[7866]<=8'd101;
		data_a[7867]<=8'd105;
		data_a[7868]<=8'd99;
		data_a[7869]<=8'd108;
		data_a[7870]<=8'd115;
		data_a[7871]<=8'd182;
		data_a[7872]<=8'd192;
		data_a[7873]<=8'd205;
		data_a[7874]<=8'd207;
		data_a[7875]<=8'd203;
		data_a[7876]<=8'd208;
		data_a[7877]<=8'd84;
		data_a[7878]<=8'd56;
		data_a[7879]<=8'd64;
		data_a[7880]<=8'd70;
		data_a[7881]<=8'd106;
		data_a[7882]<=8'd130;
		data_a[7883]<=8'd136;
		data_a[7884]<=8'd146;
		data_a[7885]<=8'd152;
		data_a[7886]<=8'd158;
		data_a[7887]<=8'd164;
		data_a[7888]<=8'd165;
		data_a[7889]<=8'd164;
		data_a[7890]<=8'd165;
		data_a[7891]<=8'd167;
		data_a[7892]<=8'd168;
		data_a[7893]<=8'd169;
		data_a[7894]<=8'd172;
		data_a[7895]<=8'd175;
		data_a[7896]<=8'd175;
		data_a[7897]<=8'd175;
		data_a[7898]<=8'd173;
		data_a[7899]<=8'd172;
		data_a[7900]<=8'd172;
		data_a[7901]<=8'd168;
		data_a[7902]<=8'd154;
		data_a[7903]<=8'd156;
		data_a[7904]<=8'd156;
		data_a[7905]<=8'd140;
		data_a[7906]<=8'd134;
		data_a[7907]<=8'd121;
		data_a[7908]<=8'd103;
		data_a[7909]<=8'd103;
		data_a[7910]<=8'd96;
		data_a[7911]<=8'd96;
		data_a[7912]<=8'd100;
		data_a[7913]<=8'd102;
		data_a[7914]<=8'd115;
		data_a[7915]<=8'd120;
		data_a[7916]<=8'd123;
		data_a[7917]<=8'd180;
		data_a[7918]<=8'd189;
		data_a[7919]<=8'd195;
		data_a[7920]<=8'd185;
		data_a[7921]<=8'd176;
		data_a[7922]<=8'd149;
		data_a[7923]<=8'd114;
		data_a[7924]<=8'd117;
		data_a[7925]<=8'd117;
		data_a[7926]<=8'd124;
		data_a[7927]<=8'd152;
		data_a[7928]<=8'd212;
		data_a[7929]<=8'd211;
		data_a[7930]<=8'd211;
		data_a[7931]<=8'd213;
		data_a[7932]<=8'd214;
		data_a[7933]<=8'd215;
		data_a[7934]<=8'd216;
		data_a[7935]<=8'd218;
		data_a[7936]<=8'd220;
		data_a[7937]<=8'd218;
		data_a[7938]<=8'd220;
		data_a[7939]<=8'd223;
		data_a[7940]<=8'd227;
		data_a[7941]<=8'd254;
		data_a[7942]<=8'd255;
		data_a[7943]<=8'd253;
		data_a[7944]<=8'd254;
		data_a[7945]<=8'd254;
		data_a[7946]<=8'd254;
		data_a[7947]<=8'd254;
		data_a[7948]<=8'd254;
		data_a[7949]<=8'd254;
		data_a[7950]<=8'd255;
		data_a[7951]<=8'd213;
		data_a[7952]<=8'd213;
		data_a[7953]<=8'd213;
		data_a[7954]<=8'd208;
		data_a[7955]<=8'd212;
		data_a[7956]<=8'd215;
		data_a[7957]<=8'd214;
		data_a[7958]<=8'd213;
		data_a[7959]<=8'd211;
		data_a[7960]<=8'd212;
		data_a[7961]<=8'd214;
		data_a[7962]<=8'd190;
		data_a[7963]<=8'd195;
		data_a[7964]<=8'd205;
		data_a[7965]<=8'd197;
		data_a[7966]<=8'd204;
		data_a[7967]<=8'd204;
		data_a[7968]<=8'd202;
		data_a[7969]<=8'd187;
		data_a[7970]<=8'd206;
		data_a[7971]<=8'd136;
		data_a[7972]<=8'd185;
		data_a[7973]<=8'd152;
		data_a[7974]<=8'd115;
		data_a[7975]<=8'd85;
		data_a[7976]<=8'd73;
		data_a[7977]<=8'd78;
		data_a[7978]<=8'd75;
		data_a[7979]<=8'd65;
		data_a[7980]<=8'd65;
		data_a[7981]<=8'd63;
		data_a[7982]<=8'd66;
		data_a[7983]<=8'd67;
		data_a[7984]<=8'd61;
		data_a[7985]<=8'd65;
		data_a[7986]<=8'd69;
		data_a[7987]<=8'd67;
		data_a[7988]<=8'd70;
		data_a[7989]<=8'd75;
		data_a[7990]<=8'd69;
		data_a[7991]<=8'd74;
		data_a[7992]<=8'd81;
		data_a[7993]<=8'd84;
		data_a[7994]<=8'd81;
		data_a[7995]<=8'd77;
		data_a[7996]<=8'd75;
		data_a[7997]<=8'd76;
		data_a[7998]<=8'd73;
		data_a[7999]<=8'd76;
		data_a[8000]<=8'd73;
		data_a[8001]<=8'd75;
		data_a[8002]<=8'd77;
		data_a[8003]<=8'd79;
		data_a[8004]<=8'd73;
		data_a[8005]<=8'd73;
		data_a[8006]<=8'd69;
		data_a[8007]<=8'd67;
		data_a[8008]<=8'd67;
		data_a[8009]<=8'd64;
		data_a[8010]<=8'd72;
		data_a[8011]<=8'd70;
		data_a[8012]<=8'd72;
		data_a[8013]<=8'd71;
		data_a[8014]<=8'd78;
		data_a[8015]<=8'd82;
		data_a[8016]<=8'd84;
		data_a[8017]<=8'd81;
		data_a[8018]<=8'd96;
		data_a[8019]<=8'd94;
		data_a[8020]<=8'd104;
		data_a[8021]<=8'd107;
		data_a[8022]<=8'd160;
		data_a[8023]<=8'd189;
		data_a[8024]<=8'd211;
		data_a[8025]<=8'd216;
		data_a[8026]<=8'd201;
		data_a[8027]<=8'd67;
		data_a[8028]<=8'd68;
		data_a[8029]<=8'd67;
		data_a[8030]<=8'd67;
		data_a[8031]<=8'd106;
		data_a[8032]<=8'd134;
		data_a[8033]<=8'd143;
		data_a[8034]<=8'd148;
		data_a[8035]<=8'd151;
		data_a[8036]<=8'd157;
		data_a[8037]<=8'd161;
		data_a[8038]<=8'd167;
		data_a[8039]<=8'd164;
		data_a[8040]<=8'd164;
		data_a[8041]<=8'd167;
		data_a[8042]<=8'd169;
		data_a[8043]<=8'd168;
		data_a[8044]<=8'd170;
		data_a[8045]<=8'd173;
		data_a[8046]<=8'd171;
		data_a[8047]<=8'd169;
		data_a[8048]<=8'd168;
		data_a[8049]<=8'd167;
		data_a[8050]<=8'd165;
		data_a[8051]<=8'd163;
		data_a[8052]<=8'd146;
		data_a[8053]<=8'd146;
		data_a[8054]<=8'd142;
		data_a[8055]<=8'd124;
		data_a[8056]<=8'd112;
		data_a[8057]<=8'd106;
		data_a[8058]<=8'd79;
		data_a[8059]<=8'd84;
		data_a[8060]<=8'd76;
		data_a[8061]<=8'd77;
		data_a[8062]<=8'd81;
		data_a[8063]<=8'd89;
		data_a[8064]<=8'd97;
		data_a[8065]<=8'd99;
		data_a[8066]<=8'd105;
		data_a[8067]<=8'd108;
		data_a[8068]<=8'd162;
		data_a[8069]<=8'd194;
		data_a[8070]<=8'd187;
		data_a[8071]<=8'd181;
		data_a[8072]<=8'd163;
		data_a[8073]<=8'd125;
		data_a[8074]<=8'd115;
		data_a[8075]<=8'd116;
		data_a[8076]<=8'd119;
		data_a[8077]<=8'd140;
		data_a[8078]<=8'd211;
		data_a[8079]<=8'd211;
		data_a[8080]<=8'd211;
		data_a[8081]<=8'd213;
		data_a[8082]<=8'd214;
		data_a[8083]<=8'd214;
		data_a[8084]<=8'd216;
		data_a[8085]<=8'd217;
		data_a[8086]<=8'd218;
		data_a[8087]<=8'd220;
		data_a[8088]<=8'd217;
		data_a[8089]<=8'd226;
		data_a[8090]<=8'd221;
		data_a[8091]<=8'd247;
		data_a[8092]<=8'd255;
		data_a[8093]<=8'd254;
		data_a[8094]<=8'd255;
		data_a[8095]<=8'd255;
		data_a[8096]<=8'd255;
		data_a[8097]<=8'd255;
		data_a[8098]<=8'd255;
		data_a[8099]<=8'd255;
		data_a[8100]<=8'd255;
		data_a[8101]<=8'd214;
		data_a[8102]<=8'd212;
		data_a[8103]<=8'd213;
		data_a[8104]<=8'd214;
		data_a[8105]<=8'd217;
		data_a[8106]<=8'd214;
		data_a[8107]<=8'd211;
		data_a[8108]<=8'd211;
		data_a[8109]<=8'd210;
		data_a[8110]<=8'd205;
		data_a[8111]<=8'd205;
		data_a[8112]<=8'd208;
		data_a[8113]<=8'd211;
		data_a[8114]<=8'd180;
		data_a[8115]<=8'd209;
		data_a[8116]<=8'd203;
		data_a[8117]<=8'd201;
		data_a[8118]<=8'd208;
		data_a[8119]<=8'd187;
		data_a[8120]<=8'd188;
		data_a[8121]<=8'd167;
		data_a[8122]<=8'd124;
		data_a[8123]<=8'd139;
		data_a[8124]<=8'd140;
		data_a[8125]<=8'd85;
		data_a[8126]<=8'd75;
		data_a[8127]<=8'd68;
		data_a[8128]<=8'd69;
		data_a[8129]<=8'd69;
		data_a[8130]<=8'd69;
		data_a[8131]<=8'd67;
		data_a[8132]<=8'd64;
		data_a[8133]<=8'd59;
		data_a[8134]<=8'd73;
		data_a[8135]<=8'd77;
		data_a[8136]<=8'd73;
		data_a[8137]<=8'd75;
		data_a[8138]<=8'd74;
		data_a[8139]<=8'd76;
		data_a[8140]<=8'd77;
		data_a[8141]<=8'd83;
		data_a[8142]<=8'd91;
		data_a[8143]<=8'd94;
		data_a[8144]<=8'd91;
		data_a[8145]<=8'd85;
		data_a[8146]<=8'd82;
		data_a[8147]<=8'd80;
		data_a[8148]<=8'd78;
		data_a[8149]<=8'd79;
		data_a[8150]<=8'd79;
		data_a[8151]<=8'd82;
		data_a[8152]<=8'd78;
		data_a[8153]<=8'd81;
		data_a[8154]<=8'd77;
		data_a[8155]<=8'd73;
		data_a[8156]<=8'd74;
		data_a[8157]<=8'd74;
		data_a[8158]<=8'd72;
		data_a[8159]<=8'd70;
		data_a[8160]<=8'd73;
		data_a[8161]<=8'd72;
		data_a[8162]<=8'd72;
		data_a[8163]<=8'd72;
		data_a[8164]<=8'd69;
		data_a[8165]<=8'd65;
		data_a[8166]<=8'd76;
		data_a[8167]<=8'd81;
		data_a[8168]<=8'd77;
		data_a[8169]<=8'd88;
		data_a[8170]<=8'd107;
		data_a[8171]<=8'd91;
		data_a[8172]<=8'd101;
		data_a[8173]<=8'd146;
		data_a[8174]<=8'd196;
		data_a[8175]<=8'd204;
		data_a[8176]<=8'd210;
		data_a[8177]<=8'd68;
		data_a[8178]<=8'd63;
		data_a[8179]<=8'd63;
		data_a[8180]<=8'd71;
		data_a[8181]<=8'd106;
		data_a[8182]<=8'd130;
		data_a[8183]<=8'd139;
		data_a[8184]<=8'd142;
		data_a[8185]<=8'd148;
		data_a[8186]<=8'd160;
		data_a[8187]<=8'd163;
		data_a[8188]<=8'd166;
		data_a[8189]<=8'd165;
		data_a[8190]<=8'd164;
		data_a[8191]<=8'd164;
		data_a[8192]<=8'd165;
		data_a[8193]<=8'd165;
		data_a[8194]<=8'd165;
		data_a[8195]<=8'd165;
		data_a[8196]<=8'd167;
		data_a[8197]<=8'd168;
		data_a[8198]<=8'd166;
		data_a[8199]<=8'd163;
		data_a[8200]<=8'd161;
		data_a[8201]<=8'd159;
		data_a[8202]<=8'd148;
		data_a[8203]<=8'd139;
		data_a[8204]<=8'd130;
		data_a[8205]<=8'd113;
		data_a[8206]<=8'd89;
		data_a[8207]<=8'd97;
		data_a[8208]<=8'd81;
		data_a[8209]<=8'd87;
		data_a[8210]<=8'd83;
		data_a[8211]<=8'd80;
		data_a[8212]<=8'd81;
		data_a[8213]<=8'd92;
		data_a[8214]<=8'd99;
		data_a[8215]<=8'd103;
		data_a[8216]<=8'd101;
		data_a[8217]<=8'd116;
		data_a[8218]<=8'd104;
		data_a[8219]<=8'd155;
		data_a[8220]<=8'd194;
		data_a[8221]<=8'd189;
		data_a[8222]<=8'd175;
		data_a[8223]<=8'd144;
		data_a[8224]<=8'd112;
		data_a[8225]<=8'd113;
		data_a[8226]<=8'd119;
		data_a[8227]<=8'd128;
		data_a[8228]<=8'd205;
		data_a[8229]<=8'd210;
		data_a[8230]<=8'd214;
		data_a[8231]<=8'd212;
		data_a[8232]<=8'd212;
		data_a[8233]<=8'd215;
		data_a[8234]<=8'd216;
		data_a[8235]<=8'd215;
		data_a[8236]<=8'd218;
		data_a[8237]<=8'd217;
		data_a[8238]<=8'd223;
		data_a[8239]<=8'd218;
		data_a[8240]<=8'd223;
		data_a[8241]<=8'd227;
		data_a[8242]<=8'd255;
		data_a[8243]<=8'd255;
		data_a[8244]<=8'd253;
		data_a[8245]<=8'd255;
		data_a[8246]<=8'd255;
		data_a[8247]<=8'd255;
		data_a[8248]<=8'd255;
		data_a[8249]<=8'd254;
		data_a[8250]<=8'd253;
		data_a[8251]<=8'd217;
		data_a[8252]<=8'd215;
		data_a[8253]<=8'd214;
		data_a[8254]<=8'd216;
		data_a[8255]<=8'd217;
		data_a[8256]<=8'd212;
		data_a[8257]<=8'd215;
		data_a[8258]<=8'd216;
		data_a[8259]<=8'd203;
		data_a[8260]<=8'd204;
		data_a[8261]<=8'd207;
		data_a[8262]<=8'd200;
		data_a[8263]<=8'd171;
		data_a[8264]<=8'd196;
		data_a[8265]<=8'd188;
		data_a[8266]<=8'd186;
		data_a[8267]<=8'd196;
		data_a[8268]<=8'd196;
		data_a[8269]<=8'd192;
		data_a[8270]<=8'd200;
		data_a[8271]<=8'd179;
		data_a[8272]<=8'd176;
		data_a[8273]<=8'd138;
		data_a[8274]<=8'd102;
		data_a[8275]<=8'd79;
		data_a[8276]<=8'd69;
		data_a[8277]<=8'd64;
		data_a[8278]<=8'd63;
		data_a[8279]<=8'd66;
		data_a[8280]<=8'd60;
		data_a[8281]<=8'd65;
		data_a[8282]<=8'd65;
		data_a[8283]<=8'd66;
		data_a[8284]<=8'd72;
		data_a[8285]<=8'd77;
		data_a[8286]<=8'd79;
		data_a[8287]<=8'd82;
		data_a[8288]<=8'd86;
		data_a[8289]<=8'd92;
		data_a[8290]<=8'd97;
		data_a[8291]<=8'd100;
		data_a[8292]<=8'd99;
		data_a[8293]<=8'd95;
		data_a[8294]<=8'd94;
		data_a[8295]<=8'd97;
		data_a[8296]<=8'd96;
		data_a[8297]<=8'd90;
		data_a[8298]<=8'd90;
		data_a[8299]<=8'd88;
		data_a[8300]<=8'd91;
		data_a[8301]<=8'd97;
		data_a[8302]<=8'd86;
		data_a[8303]<=8'd90;
		data_a[8304]<=8'd89;
		data_a[8305]<=8'd81;
		data_a[8306]<=8'd78;
		data_a[8307]<=8'd80;
		data_a[8308]<=8'd75;
		data_a[8309]<=8'd75;
		data_a[8310]<=8'd71;
		data_a[8311]<=8'd71;
		data_a[8312]<=8'd67;
		data_a[8313]<=8'd69;
		data_a[8314]<=8'd69;
		data_a[8315]<=8'd70;
		data_a[8316]<=8'd71;
		data_a[8317]<=8'd75;
		data_a[8318]<=8'd89;
		data_a[8319]<=8'd82;
		data_a[8320]<=8'd92;
		data_a[8321]<=8'd97;
		data_a[8322]<=8'd89;
		data_a[8323]<=8'd118;
		data_a[8324]<=8'd201;
		data_a[8325]<=8'd200;
		data_a[8326]<=8'd199;
		data_a[8327]<=8'd66;
		data_a[8328]<=8'd67;
		data_a[8329]<=8'd66;
		data_a[8330]<=8'd73;
		data_a[8331]<=8'd104;
		data_a[8332]<=8'd128;
		data_a[8333]<=8'd140;
		data_a[8334]<=8'd142;
		data_a[8335]<=8'd149;
		data_a[8336]<=8'd158;
		data_a[8337]<=8'd157;
		data_a[8338]<=8'd163;
		data_a[8339]<=8'd164;
		data_a[8340]<=8'd162;
		data_a[8341]<=8'd159;
		data_a[8342]<=8'd158;
		data_a[8343]<=8'd159;
		data_a[8344]<=8'd157;
		data_a[8345]<=8'd155;
		data_a[8346]<=8'd161;
		data_a[8347]<=8'd164;
		data_a[8348]<=8'd161;
		data_a[8349]<=8'd155;
		data_a[8350]<=8'd156;
		data_a[8351]<=8'd151;
		data_a[8352]<=8'd148;
		data_a[8353]<=8'd129;
		data_a[8354]<=8'd109;
		data_a[8355]<=8'd112;
		data_a[8356]<=8'd89;
		data_a[8357]<=8'd102;
		data_a[8358]<=8'd86;
		data_a[8359]<=8'd84;
		data_a[8360]<=8'd96;
		data_a[8361]<=8'd105;
		data_a[8362]<=8'd111;
		data_a[8363]<=8'd112;
		data_a[8364]<=8'd115;
		data_a[8365]<=8'd116;
		data_a[8366]<=8'd119;
		data_a[8367]<=8'd117;
		data_a[8368]<=8'd119;
		data_a[8369]<=8'd131;
		data_a[8370]<=8'd201;
		data_a[8371]<=8'd197;
		data_a[8372]<=8'd182;
		data_a[8373]<=8'd161;
		data_a[8374]<=8'd109;
		data_a[8375]<=8'd111;
		data_a[8376]<=8'd121;
		data_a[8377]<=8'd119;
		data_a[8378]<=8'd197;
		data_a[8379]<=8'd208;
		data_a[8380]<=8'd214;
		data_a[8381]<=8'd210;
		data_a[8382]<=8'd209;
		data_a[8383]<=8'd214;
		data_a[8384]<=8'd216;
		data_a[8385]<=8'd213;
		data_a[8386]<=8'd216;
		data_a[8387]<=8'd217;
		data_a[8388]<=8'd218;
		data_a[8389]<=8'd221;
		data_a[8390]<=8'd225;
		data_a[8391]<=8'd229;
		data_a[8392]<=8'd255;
		data_a[8393]<=8'd254;
		data_a[8394]<=8'd255;
		data_a[8395]<=8'd255;
		data_a[8396]<=8'd255;
		data_a[8397]<=8'd249;
		data_a[8398]<=8'd241;
		data_a[8399]<=8'd235;
		data_a[8400]<=8'd255;
		data_a[8401]<=8'd216;
		data_a[8402]<=8'd218;
		data_a[8403]<=8'd214;
		data_a[8404]<=8'd219;
		data_a[8405]<=8'd214;
		data_a[8406]<=8'd211;
		data_a[8407]<=8'd216;
		data_a[8408]<=8'd213;
		data_a[8409]<=8'd211;
		data_a[8410]<=8'd193;
		data_a[8411]<=8'd187;
		data_a[8412]<=8'd210;
		data_a[8413]<=8'd206;
		data_a[8414]<=8'd207;
		data_a[8415]<=8'd198;
		data_a[8416]<=8'd205;
		data_a[8417]<=8'd174;
		data_a[8418]<=8'd201;
		data_a[8419]<=8'd192;
		data_a[8420]<=8'd188;
		data_a[8421]<=8'd126;
		data_a[8422]<=8'd155;
		data_a[8423]<=8'd116;
		data_a[8424]<=8'd87;
		data_a[8425]<=8'd70;
		data_a[8426]<=8'd70;
		data_a[8427]<=8'd69;
		data_a[8428]<=8'd61;
		data_a[8429]<=8'd62;
		data_a[8430]<=8'd61;
		data_a[8431]<=8'd62;
		data_a[8432]<=8'd66;
		data_a[8433]<=8'd72;
		data_a[8434]<=8'd79;
		data_a[8435]<=8'd93;
		data_a[8436]<=8'd83;
		data_a[8437]<=8'd97;
		data_a[8438]<=8'd96;
		data_a[8439]<=8'd97;
		data_a[8440]<=8'd116;
		data_a[8441]<=8'd113;
		data_a[8442]<=8'd112;
		data_a[8443]<=8'd123;
		data_a[8444]<=8'd105;
		data_a[8445]<=8'd109;
		data_a[8446]<=8'd106;
		data_a[8447]<=8'd108;
		data_a[8448]<=8'd104;
		data_a[8449]<=8'd108;
		data_a[8450]<=8'd112;
		data_a[8451]<=8'd123;
		data_a[8452]<=8'd110;
		data_a[8453]<=8'd98;
		data_a[8454]<=8'd99;
		data_a[8455]<=8'd93;
		data_a[8456]<=8'd82;
		data_a[8457]<=8'd87;
		data_a[8458]<=8'd72;
		data_a[8459]<=8'd79;
		data_a[8460]<=8'd70;
		data_a[8461]<=8'd67;
		data_a[8462]<=8'd70;
		data_a[8463]<=8'd70;
		data_a[8464]<=8'd69;
		data_a[8465]<=8'd70;
		data_a[8466]<=8'd69;
		data_a[8467]<=8'd82;
		data_a[8468]<=8'd99;
		data_a[8469]<=8'd112;
		data_a[8470]<=8'd117;
		data_a[8471]<=8'd85;
		data_a[8472]<=8'd85;
		data_a[8473]<=8'd101;
		data_a[8474]<=8'd188;
		data_a[8475]<=8'd206;
		data_a[8476]<=8'd212;
		data_a[8477]<=8'd74;
		data_a[8478]<=8'd57;
		data_a[8479]<=8'd66;
		data_a[8480]<=8'd73;
		data_a[8481]<=8'd102;
		data_a[8482]<=8'd133;
		data_a[8483]<=8'd135;
		data_a[8484]<=8'd144;
		data_a[8485]<=8'd143;
		data_a[8486]<=8'd157;
		data_a[8487]<=8'd156;
		data_a[8488]<=8'd164;
		data_a[8489]<=8'd161;
		data_a[8490]<=8'd158;
		data_a[8491]<=8'd154;
		data_a[8492]<=8'd157;
		data_a[8493]<=8'd149;
		data_a[8494]<=8'd146;
		data_a[8495]<=8'd149;
		data_a[8496]<=8'd151;
		data_a[8497]<=8'd155;
		data_a[8498]<=8'd153;
		data_a[8499]<=8'd157;
		data_a[8500]<=8'd151;
		data_a[8501]<=8'd150;
		data_a[8502]<=8'd141;
		data_a[8503]<=8'd125;
		data_a[8504]<=8'd110;
		data_a[8505]<=8'd101;
		data_a[8506]<=8'd105;
		data_a[8507]<=8'd105;
		data_a[8508]<=8'd101;
		data_a[8509]<=8'd103;
		data_a[8510]<=8'd118;
		data_a[8511]<=8'd115;
		data_a[8512]<=8'd123;
		data_a[8513]<=8'd125;
		data_a[8514]<=8'd129;
		data_a[8515]<=8'd131;
		data_a[8516]<=8'd129;
		data_a[8517]<=8'd131;
		data_a[8518]<=8'd124;
		data_a[8519]<=8'd119;
		data_a[8520]<=8'd135;
		data_a[8521]<=8'd196;
		data_a[8522]<=8'd189;
		data_a[8523]<=8'd182;
		data_a[8524]<=8'd132;
		data_a[8525]<=8'd112;
		data_a[8526]<=8'd114;
		data_a[8527]<=8'd119;
		data_a[8528]<=8'd192;
		data_a[8529]<=8'd215;
		data_a[8530]<=8'd204;
		data_a[8531]<=8'd215;
		data_a[8532]<=8'd216;
		data_a[8533]<=8'd215;
		data_a[8534]<=8'd210;
		data_a[8535]<=8'd215;
		data_a[8536]<=8'd215;
		data_a[8537]<=8'd218;
		data_a[8538]<=8'd219;
		data_a[8539]<=8'd220;
		data_a[8540]<=8'd223;
		data_a[8541]<=8'd230;
		data_a[8542]<=8'd239;
		data_a[8543]<=8'd245;
		data_a[8544]<=8'd237;
		data_a[8545]<=8'd234;
		data_a[8546]<=8'd233;
		data_a[8547]<=8'd234;
		data_a[8548]<=8'd233;
		data_a[8549]<=8'd228;
		data_a[8550]<=8'd255;
		data_a[8551]<=8'd221;
		data_a[8552]<=8'd219;
		data_a[8553]<=8'd216;
		data_a[8554]<=8'd220;
		data_a[8555]<=8'd215;
		data_a[8556]<=8'd213;
		data_a[8557]<=8'd214;
		data_a[8558]<=8'd193;
		data_a[8559]<=8'd196;
		data_a[8560]<=8'd217;
		data_a[8561]<=8'd206;
		data_a[8562]<=8'd213;
		data_a[8563]<=8'd204;
		data_a[8564]<=8'd193;
		data_a[8565]<=8'd202;
		data_a[8566]<=8'd204;
		data_a[8567]<=8'd196;
		data_a[8568]<=8'd173;
		data_a[8569]<=8'd193;
		data_a[8570]<=8'd186;
		data_a[8571]<=8'd154;
		data_a[8572]<=8'd137;
		data_a[8573]<=8'd97;
		data_a[8574]<=8'd87;
		data_a[8575]<=8'd77;
		data_a[8576]<=8'd74;
		data_a[8577]<=8'd64;
		data_a[8578]<=8'd58;
		data_a[8579]<=8'd66;
		data_a[8580]<=8'd68;
		data_a[8581]<=8'd62;
		data_a[8582]<=8'd74;
		data_a[8583]<=8'd74;
		data_a[8584]<=8'd90;
		data_a[8585]<=8'd102;
		data_a[8586]<=8'd107;
		data_a[8587]<=8'd115;
		data_a[8588]<=8'd111;
		data_a[8589]<=8'd128;
		data_a[8590]<=8'd126;
		data_a[8591]<=8'd128;
		data_a[8592]<=8'd140;
		data_a[8593]<=8'd124;
		data_a[8594]<=8'd120;
		data_a[8595]<=8'd113;
		data_a[8596]<=8'd126;
		data_a[8597]<=8'd121;
		data_a[8598]<=8'd124;
		data_a[8599]<=8'd125;
		data_a[8600]<=8'd134;
		data_a[8601]<=8'd128;
		data_a[8602]<=8'd136;
		data_a[8603]<=8'd124;
		data_a[8604]<=8'd125;
		data_a[8605]<=8'd112;
		data_a[8606]<=8'd105;
		data_a[8607]<=8'd97;
		data_a[8608]<=8'd80;
		data_a[8609]<=8'd73;
		data_a[8610]<=8'd77;
		data_a[8611]<=8'd72;
		data_a[8612]<=8'd69;
		data_a[8613]<=8'd68;
		data_a[8614]<=8'd67;
		data_a[8615]<=8'd69;
		data_a[8616]<=8'd87;
		data_a[8617]<=8'd86;
		data_a[8618]<=8'd107;
		data_a[8619]<=8'd115;
		data_a[8620]<=8'd110;
		data_a[8621]<=8'd146;
		data_a[8622]<=8'd87;
		data_a[8623]<=8'd86;
		data_a[8624]<=8'd176;
		data_a[8625]<=8'd201;
		data_a[8626]<=8'd196;
		data_a[8627]<=8'd70;
		data_a[8628]<=8'd67;
		data_a[8629]<=8'd65;
		data_a[8630]<=8'd75;
		data_a[8631]<=8'd93;
		data_a[8632]<=8'd130;
		data_a[8633]<=8'd137;
		data_a[8634]<=8'd142;
		data_a[8635]<=8'd147;
		data_a[8636]<=8'd147;
		data_a[8637]<=8'd162;
		data_a[8638]<=8'd159;
		data_a[8639]<=8'd162;
		data_a[8640]<=8'd154;
		data_a[8641]<=8'd156;
		data_a[8642]<=8'd140;
		data_a[8643]<=8'd141;
		data_a[8644]<=8'd135;
		data_a[8645]<=8'd143;
		data_a[8646]<=8'd145;
		data_a[8647]<=8'd146;
		data_a[8648]<=8'd146;
		data_a[8649]<=8'd152;
		data_a[8650]<=8'd153;
		data_a[8651]<=8'd147;
		data_a[8652]<=8'd142;
		data_a[8653]<=8'd132;
		data_a[8654]<=8'd119;
		data_a[8655]<=8'd109;
		data_a[8656]<=8'd115;
		data_a[8657]<=8'd109;
		data_a[8658]<=8'd116;
		data_a[8659]<=8'd113;
		data_a[8660]<=8'd103;
		data_a[8661]<=8'd114;
		data_a[8662]<=8'd114;
		data_a[8663]<=8'd123;
		data_a[8664]<=8'd128;
		data_a[8665]<=8'd128;
		data_a[8666]<=8'd129;
		data_a[8667]<=8'd141;
		data_a[8668]<=8'd133;
		data_a[8669]<=8'd139;
		data_a[8670]<=8'd153;
		data_a[8671]<=8'd191;
		data_a[8672]<=8'd192;
		data_a[8673]<=8'd188;
		data_a[8674]<=8'd149;
		data_a[8675]<=8'd106;
		data_a[8676]<=8'd113;
		data_a[8677]<=8'd118;
		data_a[8678]<=8'd178;
		data_a[8679]<=8'd211;
		data_a[8680]<=8'd213;
		data_a[8681]<=8'd213;
		data_a[8682]<=8'd210;
		data_a[8683]<=8'd212;
		data_a[8684]<=8'd213;
		data_a[8685]<=8'd215;
		data_a[8686]<=8'd214;
		data_a[8687]<=8'd216;
		data_a[8688]<=8'd217;
		data_a[8689]<=8'd217;
		data_a[8690]<=8'd219;
		data_a[8691]<=8'd224;
		data_a[8692]<=8'd229;
		data_a[8693]<=8'd232;
		data_a[8694]<=8'd233;
		data_a[8695]<=8'd229;
		data_a[8696]<=8'd228;
		data_a[8697]<=8'd231;
		data_a[8698]<=8'd231;
		data_a[8699]<=8'd228;
		data_a[8700]<=8'd251;
		data_a[8701]<=8'd219;
		data_a[8702]<=8'd217;
		data_a[8703]<=8'd222;
		data_a[8704]<=8'd220;
		data_a[8705]<=8'd203;
		data_a[8706]<=8'd207;
		data_a[8707]<=8'd219;
		data_a[8708]<=8'd214;
		data_a[8709]<=8'd210;
		data_a[8710]<=8'd214;
		data_a[8711]<=8'd198;
		data_a[8712]<=8'd206;
		data_a[8713]<=8'd207;
		data_a[8714]<=8'd204;
		data_a[8715]<=8'd203;
		data_a[8716]<=8'd198;
		data_a[8717]<=8'd202;
		data_a[8718]<=8'd195;
		data_a[8719]<=8'd186;
		data_a[8720]<=8'd178;
		data_a[8721]<=8'd150;
		data_a[8722]<=8'd114;
		data_a[8723]<=8'd88;
		data_a[8724]<=8'd87;
		data_a[8725]<=8'd78;
		data_a[8726]<=8'd71;
		data_a[8727]<=8'd65;
		data_a[8728]<=8'd61;
		data_a[8729]<=8'd65;
		data_a[8730]<=8'd68;
		data_a[8731]<=8'd68;
		data_a[8732]<=8'd76;
		data_a[8733]<=8'd92;
		data_a[8734]<=8'd101;
		data_a[8735]<=8'd92;
		data_a[8736]<=8'd114;
		data_a[8737]<=8'd136;
		data_a[8738]<=8'd140;
		data_a[8739]<=8'd145;
		data_a[8740]<=8'd146;
		data_a[8741]<=8'd144;
		data_a[8742]<=8'd147;
		data_a[8743]<=8'd139;
		data_a[8744]<=8'd140;
		data_a[8745]<=8'd134;
		data_a[8746]<=8'd138;
		data_a[8747]<=8'd135;
		data_a[8748]<=8'd143;
		data_a[8749]<=8'd149;
		data_a[8750]<=8'd141;
		data_a[8751]<=8'd141;
		data_a[8752]<=8'd146;
		data_a[8753]<=8'd148;
		data_a[8754]<=8'd149;
		data_a[8755]<=8'd142;
		data_a[8756]<=8'd134;
		data_a[8757]<=8'd115;
		data_a[8758]<=8'd93;
		data_a[8759]<=8'd78;
		data_a[8760]<=8'd79;
		data_a[8761]<=8'd73;
		data_a[8762]<=8'd62;
		data_a[8763]<=8'd64;
		data_a[8764]<=8'd66;
		data_a[8765]<=8'd76;
		data_a[8766]<=8'd77;
		data_a[8767]<=8'd86;
		data_a[8768]<=8'd100;
		data_a[8769]<=8'd105;
		data_a[8770]<=8'd123;
		data_a[8771]<=8'd122;
		data_a[8772]<=8'd72;
		data_a[8773]<=8'd78;
		data_a[8774]<=8'd178;
		data_a[8775]<=8'd195;
		data_a[8776]<=8'd209;
		data_a[8777]<=8'd85;
		data_a[8778]<=8'd58;
		data_a[8779]<=8'd67;
		data_a[8780]<=8'd74;
		data_a[8781]<=8'd89;
		data_a[8782]<=8'd129;
		data_a[8783]<=8'd135;
		data_a[8784]<=8'd144;
		data_a[8785]<=8'd153;
		data_a[8786]<=8'd148;
		data_a[8787]<=8'd158;
		data_a[8788]<=8'd157;
		data_a[8789]<=8'd149;
		data_a[8790]<=8'd141;
		data_a[8791]<=8'd134;
		data_a[8792]<=8'd129;
		data_a[8793]<=8'd120;
		data_a[8794]<=8'd124;
		data_a[8795]<=8'd133;
		data_a[8796]<=8'd136;
		data_a[8797]<=8'd140;
		data_a[8798]<=8'd144;
		data_a[8799]<=8'd145;
		data_a[8800]<=8'd152;
		data_a[8801]<=8'd144;
		data_a[8802]<=8'd140;
		data_a[8803]<=8'd132;
		data_a[8804]<=8'd125;
		data_a[8805]<=8'd110;
		data_a[8806]<=8'd107;
		data_a[8807]<=8'd115;
		data_a[8808]<=8'd115;
		data_a[8809]<=8'd107;
		data_a[8810]<=8'd113;
		data_a[8811]<=8'd117;
		data_a[8812]<=8'd127;
		data_a[8813]<=8'd129;
		data_a[8814]<=8'd134;
		data_a[8815]<=8'd128;
		data_a[8816]<=8'd132;
		data_a[8817]<=8'd130;
		data_a[8818]<=8'd144;
		data_a[8819]<=8'd142;
		data_a[8820]<=8'd150;
		data_a[8821]<=8'd180;
		data_a[8822]<=8'd195;
		data_a[8823]<=8'd191;
		data_a[8824]<=8'd168;
		data_a[8825]<=8'd115;
		data_a[8826]<=8'd120;
		data_a[8827]<=8'd114;
		data_a[8828]<=8'd173;
		data_a[8829]<=8'd204;
		data_a[8830]<=8'd208;
		data_a[8831]<=8'd211;
		data_a[8832]<=8'd215;
		data_a[8833]<=8'd213;
		data_a[8834]<=8'd211;
		data_a[8835]<=8'd209;
		data_a[8836]<=8'd215;
		data_a[8837]<=8'd217;
		data_a[8838]<=8'd218;
		data_a[8839]<=8'd219;
		data_a[8840]<=8'd221;
		data_a[8841]<=8'd224;
		data_a[8842]<=8'd227;
		data_a[8843]<=8'd228;
		data_a[8844]<=8'd231;
		data_a[8845]<=8'd227;
		data_a[8846]<=8'd225;
		data_a[8847]<=8'd228;
		data_a[8848]<=8'd229;
		data_a[8849]<=8'd226;
		data_a[8850]<=8'd255;
		data_a[8851]<=8'd218;
		data_a[8852]<=8'd203;
		data_a[8853]<=8'd216;
		data_a[8854]<=8'd230;
		data_a[8855]<=8'd221;
		data_a[8856]<=8'd219;
		data_a[8857]<=8'd216;
		data_a[8858]<=8'd216;
		data_a[8859]<=8'd210;
		data_a[8860]<=8'd208;
		data_a[8861]<=8'd207;
		data_a[8862]<=8'd206;
		data_a[8863]<=8'd199;
		data_a[8864]<=8'd199;
		data_a[8865]<=8'd196;
		data_a[8866]<=8'd200;
		data_a[8867]<=8'd196;
		data_a[8868]<=8'd196;
		data_a[8869]<=8'd185;
		data_a[8870]<=8'd167;
		data_a[8871]<=8'd159;
		data_a[8872]<=8'd110;
		data_a[8873]<=8'd84;
		data_a[8874]<=8'd82;
		data_a[8875]<=8'd74;
		data_a[8876]<=8'd66;
		data_a[8877]<=8'd65;
		data_a[8878]<=8'd65;
		data_a[8879]<=8'd62;
		data_a[8880]<=8'd65;
		data_a[8881]<=8'd75;
		data_a[8882]<=8'd99;
		data_a[8883]<=8'd112;
		data_a[8884]<=8'd120;
		data_a[8885]<=8'd142;
		data_a[8886]<=8'd165;
		data_a[8887]<=8'd158;
		data_a[8888]<=8'd156;
		data_a[8889]<=8'd155;
		data_a[8890]<=8'd152;
		data_a[8891]<=8'd157;
		data_a[8892]<=8'd154;
		data_a[8893]<=8'd159;
		data_a[8894]<=8'd150;
		data_a[8895]<=8'd148;
		data_a[8896]<=8'd143;
		data_a[8897]<=8'd152;
		data_a[8898]<=8'd146;
		data_a[8899]<=8'd153;
		data_a[8900]<=8'd148;
		data_a[8901]<=8'd151;
		data_a[8902]<=8'd160;
		data_a[8903]<=8'd152;
		data_a[8904]<=8'd164;
		data_a[8905]<=8'd156;
		data_a[8906]<=8'd164;
		data_a[8907]<=8'd151;
		data_a[8908]<=8'd122;
		data_a[8909]<=8'd98;
		data_a[8910]<=8'd76;
		data_a[8911]<=8'd76;
		data_a[8912]<=8'd67;
		data_a[8913]<=8'd71;
		data_a[8914]<=8'd73;
		data_a[8915]<=8'd64;
		data_a[8916]<=8'd76;
		data_a[8917]<=8'd90;
		data_a[8918]<=8'd100;
		data_a[8919]<=8'd93;
		data_a[8920]<=8'd99;
		data_a[8921]<=8'd124;
		data_a[8922]<=8'd90;
		data_a[8923]<=8'd86;
		data_a[8924]<=8'd188;
		data_a[8925]<=8'd198;
		data_a[8926]<=8'd207;
		data_a[8927]<=8'd136;
		data_a[8928]<=8'd71;
		data_a[8929]<=8'd66;
		data_a[8930]<=8'd66;
		data_a[8931]<=8'd87;
		data_a[8932]<=8'd136;
		data_a[8933]<=8'd136;
		data_a[8934]<=8'd142;
		data_a[8935]<=8'd145;
		data_a[8936]<=8'd159;
		data_a[8937]<=8'd162;
		data_a[8938]<=8'd152;
		data_a[8939]<=8'd131;
		data_a[8940]<=8'd104;
		data_a[8941]<=8'd84;
		data_a[8942]<=8'd108;
		data_a[8943]<=8'd88;
		data_a[8944]<=8'd95;
		data_a[8945]<=8'd120;
		data_a[8946]<=8'd120;
		data_a[8947]<=8'd134;
		data_a[8948]<=8'd142;
		data_a[8949]<=8'd142;
		data_a[8950]<=8'd148;
		data_a[8951]<=8'd145;
		data_a[8952]<=8'd138;
		data_a[8953]<=8'd129;
		data_a[8954]<=8'd118;
		data_a[8955]<=8'd116;
		data_a[8956]<=8'd115;
		data_a[8957]<=8'd114;
		data_a[8958]<=8'd108;
		data_a[8959]<=8'd106;
		data_a[8960]<=8'd116;
		data_a[8961]<=8'd122;
		data_a[8962]<=8'd141;
		data_a[8963]<=8'd138;
		data_a[8964]<=8'd143;
		data_a[8965]<=8'd131;
		data_a[8966]<=8'd122;
		data_a[8967]<=8'd137;
		data_a[8968]<=8'd135;
		data_a[8969]<=8'd138;
		data_a[8970]<=8'd156;
		data_a[8971]<=8'd172;
		data_a[8972]<=8'd194;
		data_a[8973]<=8'd199;
		data_a[8974]<=8'd187;
		data_a[8975]<=8'd116;
		data_a[8976]<=8'd112;
		data_a[8977]<=8'd118;
		data_a[8978]<=8'd160;
		data_a[8979]<=8'd208;
		data_a[8980]<=8'd205;
		data_a[8981]<=8'd205;
		data_a[8982]<=8'd209;
		data_a[8983]<=8'd208;
		data_a[8984]<=8'd214;
		data_a[8985]<=8'd217;
		data_a[8986]<=8'd213;
		data_a[8987]<=8'd215;
		data_a[8988]<=8'd217;
		data_a[8989]<=8'd219;
		data_a[8990]<=8'd221;
		data_a[8991]<=8'd223;
		data_a[8992]<=8'd225;
		data_a[8993]<=8'd225;
		data_a[8994]<=8'd229;
		data_a[8995]<=8'd226;
		data_a[8996]<=8'd224;
		data_a[8997]<=8'd225;
		data_a[8998]<=8'd226;
		data_a[8999]<=8'd224;
		data_a[9000]<=8'd255;
		data_a[9001]<=8'd252;
		data_a[9002]<=8'd254;
		data_a[9003]<=8'd255;
		data_a[9004]<=8'd254;
		data_a[9005]<=8'd242;
		data_a[9006]<=8'd232;
		data_a[9007]<=8'd216;
		data_a[9008]<=8'd219;
		data_a[9009]<=8'd213;
		data_a[9010]<=8'd212;
		data_a[9011]<=8'd209;
		data_a[9012]<=8'd203;
		data_a[9013]<=8'd210;
		data_a[9014]<=8'd202;
		data_a[9015]<=8'd201;
		data_a[9016]<=8'd195;
		data_a[9017]<=8'd201;
		data_a[9018]<=8'd191;
		data_a[9019]<=8'd190;
		data_a[9020]<=8'd142;
		data_a[9021]<=8'd129;
		data_a[9022]<=8'd91;
		data_a[9023]<=8'd74;
		data_a[9024]<=8'd77;
		data_a[9025]<=8'd74;
		data_a[9026]<=8'd67;
		data_a[9027]<=8'd62;
		data_a[9028]<=8'd63;
		data_a[9029]<=8'd62;
		data_a[9030]<=8'd66;
		data_a[9031]<=8'd83;
		data_a[9032]<=8'd123;
		data_a[9033]<=8'd138;
		data_a[9034]<=8'd142;
		data_a[9035]<=8'd155;
		data_a[9036]<=8'd165;
		data_a[9037]<=8'd167;
		data_a[9038]<=8'd166;
		data_a[9039]<=8'd156;
		data_a[9040]<=8'd163;
		data_a[9041]<=8'd163;
		data_a[9042]<=8'd158;
		data_a[9043]<=8'd158;
		data_a[9044]<=8'd163;
		data_a[9045]<=8'd161;
		data_a[9046]<=8'd153;
		data_a[9047]<=8'd152;
		data_a[9048]<=8'd154;
		data_a[9049]<=8'd154;
		data_a[9050]<=8'd153;
		data_a[9051]<=8'd156;
		data_a[9052]<=8'd155;
		data_a[9053]<=8'd161;
		data_a[9054]<=8'd171;
		data_a[9055]<=8'd168;
		data_a[9056]<=8'd171;
		data_a[9057]<=8'd175;
		data_a[9058]<=8'd160;
		data_a[9059]<=8'd136;
		data_a[9060]<=8'd93;
		data_a[9061]<=8'd79;
		data_a[9062]<=8'd73;
		data_a[9063]<=8'd68;
		data_a[9064]<=8'd71;
		data_a[9065]<=8'd79;
		data_a[9066]<=8'd76;
		data_a[9067]<=8'd80;
		data_a[9068]<=8'd87;
		data_a[9069]<=8'd91;
		data_a[9070]<=8'd119;
		data_a[9071]<=8'd131;
		data_a[9072]<=8'd83;
		data_a[9073]<=8'd77;
		data_a[9074]<=8'd190;
		data_a[9075]<=8'd193;
		data_a[9076]<=8'd205;
		data_a[9077]<=8'd204;
		data_a[9078]<=8'd75;
		data_a[9079]<=8'd67;
		data_a[9080]<=8'd76;
		data_a[9081]<=8'd80;
		data_a[9082]<=8'd123;
		data_a[9083]<=8'd129;
		data_a[9084]<=8'd147;
		data_a[9085]<=8'd156;
		data_a[9086]<=8'd164;
		data_a[9087]<=8'd146;
		data_a[9088]<=8'd126;
		data_a[9089]<=8'd94;
		data_a[9090]<=8'd78;
		data_a[9091]<=8'd82;
		data_a[9092]<=8'd81;
		data_a[9093]<=8'd83;
		data_a[9094]<=8'd97;
		data_a[9095]<=8'd108;
		data_a[9096]<=8'd108;
		data_a[9097]<=8'd127;
		data_a[9098]<=8'd137;
		data_a[9099]<=8'd141;
		data_a[9100]<=8'd144;
		data_a[9101]<=8'd147;
		data_a[9102]<=8'd137;
		data_a[9103]<=8'd129;
		data_a[9104]<=8'd121;
		data_a[9105]<=8'd116;
		data_a[9106]<=8'd103;
		data_a[9107]<=8'd113;
		data_a[9108]<=8'd108;
		data_a[9109]<=8'd111;
		data_a[9110]<=8'd125;
		data_a[9111]<=8'd92;
		data_a[9112]<=8'd110;
		data_a[9113]<=8'd111;
		data_a[9114]<=8'd110;
		data_a[9115]<=8'd111;
		data_a[9116]<=8'd138;
		data_a[9117]<=8'd130;
		data_a[9118]<=8'd137;
		data_a[9119]<=8'd139;
		data_a[9120]<=8'd150;
		data_a[9121]<=8'd163;
		data_a[9122]<=8'd190;
		data_a[9123]<=8'd192;
		data_a[9124]<=8'd198;
		data_a[9125]<=8'd128;
		data_a[9126]<=8'd114;
		data_a[9127]<=8'd129;
		data_a[9128]<=8'd125;
		data_a[9129]<=8'd210;
		data_a[9130]<=8'd210;
		data_a[9131]<=8'd211;
		data_a[9132]<=8'd216;
		data_a[9133]<=8'd216;
		data_a[9134]<=8'd215;
		data_a[9135]<=8'd208;
		data_a[9136]<=8'd214;
		data_a[9137]<=8'd215;
		data_a[9138]<=8'd217;
		data_a[9139]<=8'd219;
		data_a[9140]<=8'd220;
		data_a[9141]<=8'd220;
		data_a[9142]<=8'd222;
		data_a[9143]<=8'd223;
		data_a[9144]<=8'd226;
		data_a[9145]<=8'd224;
		data_a[9146]<=8'd223;
		data_a[9147]<=8'd224;
		data_a[9148]<=8'd224;
		data_a[9149]<=8'd222;
		data_a[9150]<=8'd254;
		data_a[9151]<=8'd255;
		data_a[9152]<=8'd255;
		data_a[9153]<=8'd255;
		data_a[9154]<=8'd255;
		data_a[9155]<=8'd255;
		data_a[9156]<=8'd251;
		data_a[9157]<=8'd241;
		data_a[9158]<=8'd217;
		data_a[9159]<=8'd219;
		data_a[9160]<=8'd214;
		data_a[9161]<=8'd212;
		data_a[9162]<=8'd200;
		data_a[9163]<=8'd200;
		data_a[9164]<=8'd200;
		data_a[9165]<=8'd201;
		data_a[9166]<=8'd196;
		data_a[9167]<=8'd198;
		data_a[9168]<=8'd193;
		data_a[9169]<=8'd187;
		data_a[9170]<=8'd147;
		data_a[9171]<=8'd122;
		data_a[9172]<=8'd88;
		data_a[9173]<=8'd85;
		data_a[9174]<=8'd79;
		data_a[9175]<=8'd72;
		data_a[9176]<=8'd67;
		data_a[9177]<=8'd63;
		data_a[9178]<=8'd64;
		data_a[9179]<=8'd59;
		data_a[9180]<=8'd67;
		data_a[9181]<=8'd103;
		data_a[9182]<=8'd143;
		data_a[9183]<=8'd146;
		data_a[9184]<=8'd157;
		data_a[9185]<=8'd164;
		data_a[9186]<=8'd160;
		data_a[9187]<=8'd167;
		data_a[9188]<=8'd160;
		data_a[9189]<=8'd164;
		data_a[9190]<=8'd163;
		data_a[9191]<=8'd167;
		data_a[9192]<=8'd169;
		data_a[9193]<=8'd168;
		data_a[9194]<=8'd164;
		data_a[9195]<=8'd154;
		data_a[9196]<=8'd154;
		data_a[9197]<=8'd164;
		data_a[9198]<=8'd164;
		data_a[9199]<=8'd157;
		data_a[9200]<=8'd155;
		data_a[9201]<=8'd154;
		data_a[9202]<=8'd143;
		data_a[9203]<=8'd174;
		data_a[9204]<=8'd171;
		data_a[9205]<=8'd177;
		data_a[9206]<=8'd170;
		data_a[9207]<=8'd171;
		data_a[9208]<=8'd174;
		data_a[9209]<=8'd167;
		data_a[9210]<=8'd128;
		data_a[9211]<=8'd84;
		data_a[9212]<=8'd71;
		data_a[9213]<=8'd67;
		data_a[9214]<=8'd61;
		data_a[9215]<=8'd73;
		data_a[9216]<=8'd94;
		data_a[9217]<=8'd90;
		data_a[9218]<=8'd83;
		data_a[9219]<=8'd84;
		data_a[9220]<=8'd97;
		data_a[9221]<=8'd107;
		data_a[9222]<=8'd67;
		data_a[9223]<=8'd90;
		data_a[9224]<=8'd181;
		data_a[9225]<=8'd196;
		data_a[9226]<=8'd205;
		data_a[9227]<=8'd201;
		data_a[9228]<=8'd123;
		data_a[9229]<=8'd70;
		data_a[9230]<=8'd70;
		data_a[9231]<=8'd81;
		data_a[9232]<=8'd127;
		data_a[9233]<=8'd130;
		data_a[9234]<=8'd144;
		data_a[9235]<=8'd160;
		data_a[9236]<=8'd144;
		data_a[9237]<=8'd115;
		data_a[9238]<=8'd75;
		data_a[9239]<=8'd75;
		data_a[9240]<=8'd69;
		data_a[9241]<=8'd76;
		data_a[9242]<=8'd82;
		data_a[9243]<=8'd89;
		data_a[9244]<=8'd93;
		data_a[9245]<=8'd108;
		data_a[9246]<=8'd112;
		data_a[9247]<=8'd123;
		data_a[9248]<=8'd132;
		data_a[9249]<=8'd141;
		data_a[9250]<=8'd143;
		data_a[9251]<=8'd146;
		data_a[9252]<=8'd133;
		data_a[9253]<=8'd127;
		data_a[9254]<=8'd112;
		data_a[9255]<=8'd111;
		data_a[9256]<=8'd112;
		data_a[9257]<=8'd104;
		data_a[9258]<=8'd102;
		data_a[9259]<=8'd103;
		data_a[9260]<=8'd97;
		data_a[9261]<=8'd115;
		data_a[9262]<=8'd130;
		data_a[9263]<=8'd128;
		data_a[9264]<=8'd147;
		data_a[9265]<=8'd147;
		data_a[9266]<=8'd125;
		data_a[9267]<=8'd133;
		data_a[9268]<=8'd133;
		data_a[9269]<=8'd134;
		data_a[9270]<=8'd148;
		data_a[9271]<=8'd165;
		data_a[9272]<=8'd195;
		data_a[9273]<=8'd186;
		data_a[9274]<=8'd200;
		data_a[9275]<=8'd143;
		data_a[9276]<=8'd109;
		data_a[9277]<=8'd115;
		data_a[9278]<=8'd121;
		data_a[9279]<=8'd210;
		data_a[9280]<=8'd206;
		data_a[9281]<=8'd208;
		data_a[9282]<=8'd213;
		data_a[9283]<=8'd214;
		data_a[9284]<=8'd215;
		data_a[9285]<=8'd212;
		data_a[9286]<=8'd215;
		data_a[9287]<=8'd215;
		data_a[9288]<=8'd217;
		data_a[9289]<=8'd219;
		data_a[9290]<=8'd220;
		data_a[9291]<=8'd220;
		data_a[9292]<=8'd222;
		data_a[9293]<=8'd224;
		data_a[9294]<=8'd226;
		data_a[9295]<=8'd225;
		data_a[9296]<=8'd224;
		data_a[9297]<=8'd224;
		data_a[9298]<=8'd223;
		data_a[9299]<=8'd221;
		data_a[9300]<=8'd255;
		data_a[9301]<=8'd253;
		data_a[9302]<=8'd252;
		data_a[9303]<=8'd254;
		data_a[9304]<=8'd255;
		data_a[9305]<=8'd255;
		data_a[9306]<=8'd254;
		data_a[9307]<=8'd253;
		data_a[9308]<=8'd254;
		data_a[9309]<=8'd236;
		data_a[9310]<=8'd214;
		data_a[9311]<=8'd214;
		data_a[9312]<=8'd211;
		data_a[9313]<=8'd197;
		data_a[9314]<=8'd200;
		data_a[9315]<=8'd202;
		data_a[9316]<=8'd198;
		data_a[9317]<=8'd196;
		data_a[9318]<=8'd196;
		data_a[9319]<=8'd192;
		data_a[9320]<=8'd141;
		data_a[9321]<=8'd111;
		data_a[9322]<=8'd72;
		data_a[9323]<=8'd81;
		data_a[9324]<=8'd79;
		data_a[9325]<=8'd69;
		data_a[9326]<=8'd67;
		data_a[9327]<=8'd63;
		data_a[9328]<=8'd66;
		data_a[9329]<=8'd60;
		data_a[9330]<=8'd69;
		data_a[9331]<=8'd123;
		data_a[9332]<=8'd147;
		data_a[9333]<=8'd150;
		data_a[9334]<=8'd161;
		data_a[9335]<=8'd162;
		data_a[9336]<=8'd157;
		data_a[9337]<=8'd167;
		data_a[9338]<=8'd159;
		data_a[9339]<=8'd167;
		data_a[9340]<=8'd167;
		data_a[9341]<=8'd164;
		data_a[9342]<=8'd162;
		data_a[9343]<=8'd170;
		data_a[9344]<=8'd165;
		data_a[9345]<=8'd157;
		data_a[9346]<=8'd153;
		data_a[9347]<=8'd161;
		data_a[9348]<=8'd160;
		data_a[9349]<=8'd156;
		data_a[9350]<=8'd163;
		data_a[9351]<=8'd156;
		data_a[9352]<=8'd159;
		data_a[9353]<=8'd170;
		data_a[9354]<=8'd171;
		data_a[9355]<=8'd171;
		data_a[9356]<=8'd176;
		data_a[9357]<=8'd168;
		data_a[9358]<=8'd170;
		data_a[9359]<=8'd171;
		data_a[9360]<=8'd152;
		data_a[9361]<=8'd109;
		data_a[9362]<=8'd78;
		data_a[9363]<=8'd77;
		data_a[9364]<=8'd73;
		data_a[9365]<=8'd77;
		data_a[9366]<=8'd80;
		data_a[9367]<=8'd68;
		data_a[9368]<=8'd80;
		data_a[9369]<=8'd89;
		data_a[9370]<=8'd81;
		data_a[9371]<=8'd86;
		data_a[9372]<=8'd90;
		data_a[9373]<=8'd195;
		data_a[9374]<=8'd199;
		data_a[9375]<=8'd182;
		data_a[9376]<=8'd204;
		data_a[9377]<=8'd201;
		data_a[9378]<=8'd216;
		data_a[9379]<=8'd68;
		data_a[9380]<=8'd67;
		data_a[9381]<=8'd83;
		data_a[9382]<=8'd122;
		data_a[9383]<=8'd128;
		data_a[9384]<=8'd148;
		data_a[9385]<=8'd146;
		data_a[9386]<=8'd113;
		data_a[9387]<=8'd81;
		data_a[9388]<=8'd73;
		data_a[9389]<=8'd73;
		data_a[9390]<=8'd81;
		data_a[9391]<=8'd79;
		data_a[9392]<=8'd92;
		data_a[9393]<=8'd93;
		data_a[9394]<=8'd106;
		data_a[9395]<=8'd108;
		data_a[9396]<=8'd114;
		data_a[9397]<=8'd117;
		data_a[9398]<=8'd128;
		data_a[9399]<=8'd136;
		data_a[9400]<=8'd144;
		data_a[9401]<=8'd150;
		data_a[9402]<=8'd137;
		data_a[9403]<=8'd124;
		data_a[9404]<=8'd114;
		data_a[9405]<=8'd108;
		data_a[9406]<=8'd107;
		data_a[9407]<=8'd105;
		data_a[9408]<=8'd94;
		data_a[9409]<=8'd94;
		data_a[9410]<=8'd97;
		data_a[9411]<=8'd109;
		data_a[9412]<=8'd80;
		data_a[9413]<=8'd74;
		data_a[9414]<=8'd77;
		data_a[9415]<=8'd103;
		data_a[9416]<=8'd126;
		data_a[9417]<=8'd113;
		data_a[9418]<=8'd118;
		data_a[9419]<=8'd146;
		data_a[9420]<=8'd140;
		data_a[9421]<=8'd151;
		data_a[9422]<=8'd178;
		data_a[9423]<=8'd191;
		data_a[9424]<=8'd202;
		data_a[9425]<=8'd168;
		data_a[9426]<=8'd107;
		data_a[9427]<=8'd113;
		data_a[9428]<=8'd122;
		data_a[9429]<=8'd201;
		data_a[9430]<=8'd211;
		data_a[9431]<=8'd212;
		data_a[9432]<=8'd211;
		data_a[9433]<=8'd206;
		data_a[9434]<=8'd208;
		data_a[9435]<=8'd216;
		data_a[9436]<=8'd212;
		data_a[9437]<=8'd211;
		data_a[9438]<=8'd213;
		data_a[9439]<=8'd215;
		data_a[9440]<=8'd218;
		data_a[9441]<=8'd219;
		data_a[9442]<=8'd220;
		data_a[9443]<=8'd221;
		data_a[9444]<=8'd224;
		data_a[9445]<=8'd222;
		data_a[9446]<=8'd221;
		data_a[9447]<=8'd221;
		data_a[9448]<=8'd221;
		data_a[9449]<=8'd220;
		data_a[9450]<=8'd253;
		data_a[9451]<=8'd255;
		data_a[9452]<=8'd255;
		data_a[9453]<=8'd255;
		data_a[9454]<=8'd252;
		data_a[9455]<=8'd255;
		data_a[9456]<=8'd254;
		data_a[9457]<=8'd255;
		data_a[9458]<=8'd255;
		data_a[9459]<=8'd253;
		data_a[9460]<=8'd251;
		data_a[9461]<=8'd210;
		data_a[9462]<=8'd200;
		data_a[9463]<=8'd203;
		data_a[9464]<=8'd198;
		data_a[9465]<=8'd198;
		data_a[9466]<=8'd196;
		data_a[9467]<=8'd193;
		data_a[9468]<=8'd190;
		data_a[9469]<=8'd195;
		data_a[9470]<=8'd142;
		data_a[9471]<=8'd95;
		data_a[9472]<=8'd75;
		data_a[9473]<=8'd68;
		data_a[9474]<=8'd71;
		data_a[9475]<=8'd69;
		data_a[9476]<=8'd71;
		data_a[9477]<=8'd60;
		data_a[9478]<=8'd63;
		data_a[9479]<=8'd65;
		data_a[9480]<=8'd76;
		data_a[9481]<=8'd132;
		data_a[9482]<=8'd140;
		data_a[9483]<=8'd152;
		data_a[9484]<=8'd156;
		data_a[9485]<=8'd157;
		data_a[9486]<=8'd159;
		data_a[9487]<=8'd167;
		data_a[9488]<=8'd161;
		data_a[9489]<=8'd160;
		data_a[9490]<=8'd159;
		data_a[9491]<=8'd161;
		data_a[9492]<=8'd165;
		data_a[9493]<=8'd163;
		data_a[9494]<=8'd163;
		data_a[9495]<=8'd157;
		data_a[9496]<=8'd156;
		data_a[9497]<=8'd154;
		data_a[9498]<=8'd157;
		data_a[9499]<=8'd166;
		data_a[9500]<=8'd159;
		data_a[9501]<=8'd167;
		data_a[9502]<=8'd166;
		data_a[9503]<=8'd164;
		data_a[9504]<=8'd171;
		data_a[9505]<=8'd173;
		data_a[9506]<=8'd164;
		data_a[9507]<=8'd169;
		data_a[9508]<=8'd169;
		data_a[9509]<=8'd167;
		data_a[9510]<=8'd162;
		data_a[9511]<=8'd143;
		data_a[9512]<=8'd87;
		data_a[9513]<=8'd68;
		data_a[9514]<=8'd63;
		data_a[9515]<=8'd63;
		data_a[9516]<=8'd69;
		data_a[9517]<=8'd70;
		data_a[9518]<=8'd69;
		data_a[9519]<=8'd86;
		data_a[9520]<=8'd107;
		data_a[9521]<=8'd85;
		data_a[9522]<=8'd132;
		data_a[9523]<=8'd177;
		data_a[9524]<=8'd180;
		data_a[9525]<=8'd190;
		data_a[9526]<=8'd201;
		data_a[9527]<=8'd206;
		data_a[9528]<=8'd209;
		data_a[9529]<=8'd51;
		data_a[9530]<=8'd65;
		data_a[9531]<=8'd82;
		data_a[9532]<=8'd116;
		data_a[9533]<=8'd130;
		data_a[9534]<=8'd151;
		data_a[9535]<=8'd108;
		data_a[9536]<=8'd90;
		data_a[9537]<=8'd82;
		data_a[9538]<=8'd71;
		data_a[9539]<=8'd65;
		data_a[9540]<=8'd83;
		data_a[9541]<=8'd89;
		data_a[9542]<=8'd104;
		data_a[9543]<=8'd104;
		data_a[9544]<=8'd113;
		data_a[9545]<=8'd101;
		data_a[9546]<=8'd107;
		data_a[9547]<=8'd109;
		data_a[9548]<=8'd123;
		data_a[9549]<=8'd129;
		data_a[9550]<=8'd147;
		data_a[9551]<=8'd160;
		data_a[9552]<=8'd148;
		data_a[9553]<=8'd125;
		data_a[9554]<=8'd107;
		data_a[9555]<=8'd110;
		data_a[9556]<=8'd108;
		data_a[9557]<=8'd99;
		data_a[9558]<=8'd86;
		data_a[9559]<=8'd96;
		data_a[9560]<=8'd89;
		data_a[9561]<=8'd68;
		data_a[9562]<=8'd72;
		data_a[9563]<=8'd71;
		data_a[9564]<=8'd76;
		data_a[9565]<=8'd80;
		data_a[9566]<=8'd76;
		data_a[9567]<=8'd92;
		data_a[9568]<=8'd101;
		data_a[9569]<=8'd110;
		data_a[9570]<=8'd136;
		data_a[9571]<=8'd152;
		data_a[9572]<=8'd169;
		data_a[9573]<=8'd192;
		data_a[9574]<=8'd190;
		data_a[9575]<=8'd194;
		data_a[9576]<=8'd113;
		data_a[9577]<=8'd108;
		data_a[9578]<=8'd130;
		data_a[9579]<=8'd193;
		data_a[9580]<=8'd207;
		data_a[9581]<=8'd202;
		data_a[9582]<=8'd208;
		data_a[9583]<=8'd213;
		data_a[9584]<=8'd212;
		data_a[9585]<=8'd210;
		data_a[9586]<=8'd214;
		data_a[9587]<=8'd212;
		data_a[9588]<=8'd213;
		data_a[9589]<=8'd216;
		data_a[9590]<=8'd219;
		data_a[9591]<=8'd220;
		data_a[9592]<=8'd220;
		data_a[9593]<=8'd220;
		data_a[9594]<=8'd217;
		data_a[9595]<=8'd215;
		data_a[9596]<=8'd214;
		data_a[9597]<=8'd215;
		data_a[9598]<=8'd217;
		data_a[9599]<=8'd217;
		data_a[9600]<=8'd253;
		data_a[9601]<=8'd255;
		data_a[9602]<=8'd254;
		data_a[9603]<=8'd254;
		data_a[9604]<=8'd255;
		data_a[9605]<=8'd255;
		data_a[9606]<=8'd253;
		data_a[9607]<=8'd255;
		data_a[9608]<=8'd253;
		data_a[9609]<=8'd253;
		data_a[9610]<=8'd248;
		data_a[9611]<=8'd255;
		data_a[9612]<=8'd214;
		data_a[9613]<=8'd204;
		data_a[9614]<=8'd196;
		data_a[9615]<=8'd202;
		data_a[9616]<=8'd195;
		data_a[9617]<=8'd200;
		data_a[9618]<=8'd188;
		data_a[9619]<=8'd194;
		data_a[9620]<=8'd139;
		data_a[9621]<=8'd74;
		data_a[9622]<=8'd71;
		data_a[9623]<=8'd75;
		data_a[9624]<=8'd77;
		data_a[9625]<=8'd66;
		data_a[9626]<=8'd66;
		data_a[9627]<=8'd63;
		data_a[9628]<=8'd60;
		data_a[9629]<=8'd61;
		data_a[9630]<=8'd107;
		data_a[9631]<=8'd137;
		data_a[9632]<=8'd155;
		data_a[9633]<=8'd154;
		data_a[9634]<=8'd157;
		data_a[9635]<=8'd165;
		data_a[9636]<=8'd151;
		data_a[9637]<=8'd158;
		data_a[9638]<=8'd159;
		data_a[9639]<=8'd156;
		data_a[9640]<=8'd155;
		data_a[9641]<=8'd154;
		data_a[9642]<=8'd152;
		data_a[9643]<=8'd157;
		data_a[9644]<=8'd158;
		data_a[9645]<=8'd153;
		data_a[9646]<=8'd163;
		data_a[9647]<=8'd159;
		data_a[9648]<=8'd159;
		data_a[9649]<=8'd160;
		data_a[9650]<=8'd167;
		data_a[9651]<=8'd164;
		data_a[9652]<=8'd163;
		data_a[9653]<=8'd168;
		data_a[9654]<=8'd164;
		data_a[9655]<=8'd162;
		data_a[9656]<=8'd169;
		data_a[9657]<=8'd162;
		data_a[9658]<=8'd163;
		data_a[9659]<=8'd162;
		data_a[9660]<=8'd165;
		data_a[9661]<=8'd152;
		data_a[9662]<=8'd102;
		data_a[9663]<=8'd72;
		data_a[9664]<=8'd72;
		data_a[9665]<=8'd64;
		data_a[9666]<=8'd61;
		data_a[9667]<=8'd56;
		data_a[9668]<=8'd61;
		data_a[9669]<=8'd71;
		data_a[9670]<=8'd85;
		data_a[9671]<=8'd82;
		data_a[9672]<=8'd137;
		data_a[9673]<=8'd141;
		data_a[9674]<=8'd161;
		data_a[9675]<=8'd191;
		data_a[9676]<=8'd202;
		data_a[9677]<=8'd202;
		data_a[9678]<=8'd204;
		data_a[9679]<=8'd66;
		data_a[9680]<=8'd67;
		data_a[9681]<=8'd72;
		data_a[9682]<=8'd118;
		data_a[9683]<=8'd129;
		data_a[9684]<=8'd152;
		data_a[9685]<=8'd104;
		data_a[9686]<=8'd81;
		data_a[9687]<=8'd77;
		data_a[9688]<=8'd71;
		data_a[9689]<=8'd79;
		data_a[9690]<=8'd92;
		data_a[9691]<=8'd101;
		data_a[9692]<=8'd110;
		data_a[9693]<=8'd106;
		data_a[9694]<=8'd106;
		data_a[9695]<=8'd108;
		data_a[9696]<=8'd106;
		data_a[9697]<=8'd108;
		data_a[9698]<=8'd120;
		data_a[9699]<=8'd132;
		data_a[9700]<=8'd147;
		data_a[9701]<=8'd170;
		data_a[9702]<=8'd161;
		data_a[9703]<=8'd129;
		data_a[9704]<=8'd106;
		data_a[9705]<=8'd104;
		data_a[9706]<=8'd99;
		data_a[9707]<=8'd94;
		data_a[9708]<=8'd92;
		data_a[9709]<=8'd103;
		data_a[9710]<=8'd87;
		data_a[9711]<=8'd78;
		data_a[9712]<=8'd80;
		data_a[9713]<=8'd71;
		data_a[9714]<=8'd74;
		data_a[9715]<=8'd113;
		data_a[9716]<=8'd85;
		data_a[9717]<=8'd82;
		data_a[9718]<=8'd93;
		data_a[9719]<=8'd109;
		data_a[9720]<=8'd132;
		data_a[9721]<=8'd140;
		data_a[9722]<=8'd171;
		data_a[9723]<=8'd186;
		data_a[9724]<=8'd195;
		data_a[9725]<=8'd198;
		data_a[9726]<=8'd127;
		data_a[9727]<=8'd118;
		data_a[9728]<=8'd122;
		data_a[9729]<=8'd169;
		data_a[9730]<=8'd235;
		data_a[9731]<=8'd204;
		data_a[9732]<=8'd210;
		data_a[9733]<=8'd213;
		data_a[9734]<=8'd210;
		data_a[9735]<=8'd212;
		data_a[9736]<=8'd209;
		data_a[9737]<=8'd212;
		data_a[9738]<=8'd214;
		data_a[9739]<=8'd214;
		data_a[9740]<=8'd212;
		data_a[9741]<=8'd211;
		data_a[9742]<=8'd213;
		data_a[9743]<=8'd215;
		data_a[9744]<=8'd218;
		data_a[9745]<=8'd217;
		data_a[9746]<=8'd214;
		data_a[9747]<=8'd217;
		data_a[9748]<=8'd211;
		data_a[9749]<=8'd210;
		data_a[9750]<=8'd252;
		data_a[9751]<=8'd255;
		data_a[9752]<=8'd255;
		data_a[9753]<=8'd254;
		data_a[9754]<=8'd253;
		data_a[9755]<=8'd252;
		data_a[9756]<=8'd255;
		data_a[9757]<=8'd252;
		data_a[9758]<=8'd255;
		data_a[9759]<=8'd255;
		data_a[9760]<=8'd249;
		data_a[9761]<=8'd254;
		data_a[9762]<=8'd255;
		data_a[9763]<=8'd202;
		data_a[9764]<=8'd194;
		data_a[9765]<=8'd187;
		data_a[9766]<=8'd195;
		data_a[9767]<=8'd195;
		data_a[9768]<=8'd160;
		data_a[9769]<=8'd184;
		data_a[9770]<=8'd123;
		data_a[9771]<=8'd79;
		data_a[9772]<=8'd72;
		data_a[9773]<=8'd71;
		data_a[9774]<=8'd70;
		data_a[9775]<=8'd59;
		data_a[9776]<=8'd60;
		data_a[9777]<=8'd61;
		data_a[9778]<=8'd59;
		data_a[9779]<=8'd63;
		data_a[9780]<=8'd113;
		data_a[9781]<=8'd148;
		data_a[9782]<=8'd144;
		data_a[9783]<=8'd156;
		data_a[9784]<=8'd158;
		data_a[9785]<=8'd157;
		data_a[9786]<=8'd160;
		data_a[9787]<=8'd152;
		data_a[9788]<=8'd148;
		data_a[9789]<=8'd156;
		data_a[9790]<=8'd152;
		data_a[9791]<=8'd151;
		data_a[9792]<=8'd153;
		data_a[9793]<=8'd155;
		data_a[9794]<=8'd157;
		data_a[9795]<=8'd153;
		data_a[9796]<=8'd156;
		data_a[9797]<=8'd153;
		data_a[9798]<=8'd155;
		data_a[9799]<=8'd157;
		data_a[9800]<=8'd159;
		data_a[9801]<=8'd160;
		data_a[9802]<=8'd159;
		data_a[9803]<=8'd160;
		data_a[9804]<=8'd162;
		data_a[9805]<=8'd159;
		data_a[9806]<=8'd161;
		data_a[9807]<=8'd165;
		data_a[9808]<=8'd167;
		data_a[9809]<=8'd155;
		data_a[9810]<=8'd158;
		data_a[9811]<=8'd160;
		data_a[9812]<=8'd122;
		data_a[9813]<=8'd78;
		data_a[9814]<=8'd64;
		data_a[9815]<=8'd65;
		data_a[9816]<=8'd60;
		data_a[9817]<=8'd64;
		data_a[9818]<=8'd75;
		data_a[9819]<=8'd72;
		data_a[9820]<=8'd74;
		data_a[9821]<=8'd97;
		data_a[9822]<=8'd115;
		data_a[9823]<=8'd151;
		data_a[9824]<=8'd183;
		data_a[9825]<=8'd184;
		data_a[9826]<=8'd198;
		data_a[9827]<=8'd207;
		data_a[9828]<=8'd203;
		data_a[9829]<=8'd84;
		data_a[9830]<=8'd62;
		data_a[9831]<=8'd72;
		data_a[9832]<=8'd114;
		data_a[9833]<=8'd135;
		data_a[9834]<=8'd133;
		data_a[9835]<=8'd90;
		data_a[9836]<=8'd81;
		data_a[9837]<=8'd75;
		data_a[9838]<=8'd110;
		data_a[9839]<=8'd113;
		data_a[9840]<=8'd107;
		data_a[9841]<=8'd111;
		data_a[9842]<=8'd99;
		data_a[9843]<=8'd101;
		data_a[9844]<=8'd105;
		data_a[9845]<=8'd100;
		data_a[9846]<=8'd103;
		data_a[9847]<=8'd105;
		data_a[9848]<=8'd109;
		data_a[9849]<=8'd125;
		data_a[9850]<=8'd161;
		data_a[9851]<=8'd187;
		data_a[9852]<=8'd167;
		data_a[9853]<=8'd135;
		data_a[9854]<=8'd111;
		data_a[9855]<=8'd97;
		data_a[9856]<=8'd98;
		data_a[9857]<=8'd89;
		data_a[9858]<=8'd94;
		data_a[9859]<=8'd77;
		data_a[9860]<=8'd125;
		data_a[9861]<=8'd78;
		data_a[9862]<=8'd84;
		data_a[9863]<=8'd89;
		data_a[9864]<=8'd79;
		data_a[9865]<=8'd88;
		data_a[9866]<=8'd110;
		data_a[9867]<=8'd116;
		data_a[9868]<=8'd130;
		data_a[9869]<=8'd123;
		data_a[9870]<=8'd150;
		data_a[9871]<=8'd163;
		data_a[9872]<=8'd174;
		data_a[9873]<=8'd184;
		data_a[9874]<=8'd194;
		data_a[9875]<=8'd205;
		data_a[9876]<=8'd160;
		data_a[9877]<=8'd116;
		data_a[9878]<=8'd130;
		data_a[9879]<=8'd161;
		data_a[9880]<=8'd189;
		data_a[9881]<=8'd208;
		data_a[9882]<=8'd206;
		data_a[9883]<=8'd208;
		data_a[9884]<=8'd209;
		data_a[9885]<=8'd205;
		data_a[9886]<=8'd209;
		data_a[9887]<=8'd207;
		data_a[9888]<=8'd207;
		data_a[9889]<=8'd210;
		data_a[9890]<=8'd215;
		data_a[9891]<=8'd217;
		data_a[9892]<=8'd216;
		data_a[9893]<=8'd213;
		data_a[9894]<=8'd214;
		data_a[9895]<=8'd213;
		data_a[9896]<=8'd209;
		data_a[9897]<=8'd210;
		data_a[9898]<=8'd203;
		data_a[9899]<=8'd201;
		data_a[9900]<=8'd255;
		data_a[9901]<=8'd248;
		data_a[9902]<=8'd254;
		data_a[9903]<=8'd254;
		data_a[9904]<=8'd255;
		data_a[9905]<=8'd252;
		data_a[9906]<=8'd255;
		data_a[9907]<=8'd255;
		data_a[9908]<=8'd255;
		data_a[9909]<=8'd254;
		data_a[9910]<=8'd250;
		data_a[9911]<=8'd255;
		data_a[9912]<=8'd242;
		data_a[9913]<=8'd237;
		data_a[9914]<=8'd240;
		data_a[9915]<=8'd164;
		data_a[9916]<=8'd179;
		data_a[9917]<=8'd189;
		data_a[9918]<=8'd193;
		data_a[9919]<=8'd187;
		data_a[9920]<=8'd117;
		data_a[9921]<=8'd75;
		data_a[9922]<=8'd72;
		data_a[9923]<=8'd76;
		data_a[9924]<=8'd69;
		data_a[9925]<=8'd63;
		data_a[9926]<=8'd64;
		data_a[9927]<=8'd63;
		data_a[9928]<=8'd61;
		data_a[9929]<=8'd71;
		data_a[9930]<=8'd123;
		data_a[9931]<=8'd156;
		data_a[9932]<=8'd147;
		data_a[9933]<=8'd160;
		data_a[9934]<=8'd157;
		data_a[9935]<=8'd154;
		data_a[9936]<=8'd162;
		data_a[9937]<=8'd151;
		data_a[9938]<=8'd141;
		data_a[9939]<=8'd155;
		data_a[9940]<=8'd152;
		data_a[9941]<=8'd152;
		data_a[9942]<=8'd155;
		data_a[9943]<=8'd150;
		data_a[9944]<=8'd154;
		data_a[9945]<=8'd153;
		data_a[9946]<=8'd152;
		data_a[9947]<=8'd153;
		data_a[9948]<=8'd153;
		data_a[9949]<=8'd155;
		data_a[9950]<=8'd153;
		data_a[9951]<=8'd157;
		data_a[9952]<=8'd155;
		data_a[9953]<=8'd153;
		data_a[9954]<=8'd159;
		data_a[9955]<=8'd156;
		data_a[9956]<=8'd154;
		data_a[9957]<=8'd158;
		data_a[9958]<=8'd164;
		data_a[9959]<=8'd156;
		data_a[9960]<=8'd160;
		data_a[9961]<=8'd160;
		data_a[9962]<=8'd135;
		data_a[9963]<=8'd88;
		data_a[9964]<=8'd68;
		data_a[9965]<=8'd64;
		data_a[9966]<=8'd66;
		data_a[9967]<=8'd59;
		data_a[9968]<=8'd62;
		data_a[9969]<=8'd68;
		data_a[9970]<=8'd83;
		data_a[9971]<=8'd86;
		data_a[9972]<=8'd91;
		data_a[9973]<=8'd118;
		data_a[9974]<=8'd159;
		data_a[9975]<=8'd198;
		data_a[9976]<=8'd197;
		data_a[9977]<=8'd203;
		data_a[9978]<=8'd204;
		data_a[9979]<=8'd112;
		data_a[9980]<=8'd75;
		data_a[9981]<=8'd77;
		data_a[9982]<=8'd110;
		data_a[9983]<=8'd126;
		data_a[9984]<=8'd98;
		data_a[9985]<=8'd83;
		data_a[9986]<=8'd99;
		data_a[9987]<=8'd108;
		data_a[9988]<=8'd118;
		data_a[9989]<=8'd110;
		data_a[9990]<=8'd108;
		data_a[9991]<=8'd108;
		data_a[9992]<=8'd102;
		data_a[9993]<=8'd106;
		data_a[9994]<=8'd102;
		data_a[9995]<=8'd96;
		data_a[9996]<=8'd97;
		data_a[9997]<=8'd97;
		data_a[9998]<=8'd107;
		data_a[9999]<=8'd121;
		data_a[10000]<=8'd159;
		data_a[10001]<=8'd188;
		data_a[10002]<=8'd179;
		data_a[10003]<=8'd155;
		data_a[10004]<=8'd106;
		data_a[10005]<=8'd97;
		data_a[10006]<=8'd100;
		data_a[10007]<=8'd90;
		data_a[10008]<=8'd81;
		data_a[10009]<=8'd92;
		data_a[10010]<=8'd132;
		data_a[10011]<=8'd81;
		data_a[10012]<=8'd96;
		data_a[10013]<=8'd68;
		data_a[10014]<=8'd88;
		data_a[10015]<=8'd99;
		data_a[10016]<=8'd108;
		data_a[10017]<=8'd128;
		data_a[10018]<=8'd137;
		data_a[10019]<=8'd159;
		data_a[10020]<=8'd167;
		data_a[10021]<=8'd182;
		data_a[10022]<=8'd187;
		data_a[10023]<=8'd184;
		data_a[10024]<=8'd203;
		data_a[10025]<=8'd200;
		data_a[10026]<=8'd190;
		data_a[10027]<=8'd109;
		data_a[10028]<=8'd120;
		data_a[10029]<=8'd153;
		data_a[10030]<=8'd177;
		data_a[10031]<=8'd223;
		data_a[10032]<=8'd205;
		data_a[10033]<=8'd203;
		data_a[10034]<=8'd203;
		data_a[10035]<=8'd206;
		data_a[10036]<=8'd204;
		data_a[10037]<=8'd205;
		data_a[10038]<=8'd206;
		data_a[10039]<=8'd207;
		data_a[10040]<=8'd208;
		data_a[10041]<=8'd209;
		data_a[10042]<=8'd209;
		data_a[10043]<=8'd209;
		data_a[10044]<=8'd198;
		data_a[10045]<=8'd199;
		data_a[10046]<=8'd199;
		data_a[10047]<=8'd205;
		data_a[10048]<=8'd206;
		data_a[10049]<=8'd208;
		data_a[10050]<=8'd249;
		data_a[10051]<=8'd255;
		data_a[10052]<=8'd255;
		data_a[10053]<=8'd255;
		data_a[10054]<=8'd253;
		data_a[10055]<=8'd255;
		data_a[10056]<=8'd252;
		data_a[10057]<=8'd253;
		data_a[10058]<=8'd253;
		data_a[10059]<=8'd255;
		data_a[10060]<=8'd248;
		data_a[10061]<=8'd248;
		data_a[10062]<=8'd231;
		data_a[10063]<=8'd177;
		data_a[10064]<=8'd193;
		data_a[10065]<=8'd193;
		data_a[10066]<=8'd190;
		data_a[10067]<=8'd189;
		data_a[10068]<=8'd190;
		data_a[10069]<=8'd175;
		data_a[10070]<=8'd100;
		data_a[10071]<=8'd74;
		data_a[10072]<=8'd68;
		data_a[10073]<=8'd70;
		data_a[10074]<=8'd62;
		data_a[10075]<=8'd64;
		data_a[10076]<=8'd65;
		data_a[10077]<=8'd58;
		data_a[10078]<=8'd56;
		data_a[10079]<=8'd74;
		data_a[10080]<=8'd124;
		data_a[10081]<=8'd148;
		data_a[10082]<=8'd160;
		data_a[10083]<=8'd161;
		data_a[10084]<=8'd152;
		data_a[10085]<=8'd158;
		data_a[10086]<=8'd156;
		data_a[10087]<=8'd155;
		data_a[10088]<=8'd146;
		data_a[10089]<=8'd154;
		data_a[10090]<=8'd151;
		data_a[10091]<=8'd154;
		data_a[10092]<=8'd154;
		data_a[10093]<=8'd148;
		data_a[10094]<=8'd152;
		data_a[10095]<=8'd151;
		data_a[10096]<=8'd150;
		data_a[10097]<=8'd150;
		data_a[10098]<=8'd152;
		data_a[10099]<=8'd152;
		data_a[10100]<=8'd151;
		data_a[10101]<=8'd155;
		data_a[10102]<=8'd152;
		data_a[10103]<=8'd148;
		data_a[10104]<=8'd152;
		data_a[10105]<=8'd151;
		data_a[10106]<=8'd155;
		data_a[10107]<=8'd147;
		data_a[10108]<=8'd148;
		data_a[10109]<=8'd145;
		data_a[10110]<=8'd149;
		data_a[10111]<=8'd147;
		data_a[10112]<=8'd141;
		data_a[10113]<=8'd103;
		data_a[10114]<=8'd65;
		data_a[10115]<=8'd64;
		data_a[10116]<=8'd54;
		data_a[10117]<=8'd72;
		data_a[10118]<=8'd70;
		data_a[10119]<=8'd83;
		data_a[10120]<=8'd75;
		data_a[10121]<=8'd95;
		data_a[10122]<=8'd98;
		data_a[10123]<=8'd103;
		data_a[10124]<=8'd173;
		data_a[10125]<=8'd207;
		data_a[10126]<=8'd198;
		data_a[10127]<=8'd197;
		data_a[10128]<=8'd203;
		data_a[10129]<=8'd147;
		data_a[10130]<=8'd70;
		data_a[10131]<=8'd69;
		data_a[10132]<=8'd114;
		data_a[10133]<=8'd125;
		data_a[10134]<=8'd89;
		data_a[10135]<=8'd96;
		data_a[10136]<=8'd106;
		data_a[10137]<=8'd119;
		data_a[10138]<=8'd121;
		data_a[10139]<=8'd112;
		data_a[10140]<=8'd111;
		data_a[10141]<=8'd104;
		data_a[10142]<=8'd99;
		data_a[10143]<=8'd92;
		data_a[10144]<=8'd85;
		data_a[10145]<=8'd92;
		data_a[10146]<=8'd91;
		data_a[10147]<=8'd91;
		data_a[10148]<=8'd99;
		data_a[10149]<=8'd110;
		data_a[10150]<=8'd162;
		data_a[10151]<=8'd191;
		data_a[10152]<=8'd191;
		data_a[10153]<=8'd174;
		data_a[10154]<=8'd132;
		data_a[10155]<=8'd102;
		data_a[10156]<=8'd90;
		data_a[10157]<=8'd94;
		data_a[10158]<=8'd78;
		data_a[10159]<=8'd99;
		data_a[10160]<=8'd118;
		data_a[10161]<=8'd97;
		data_a[10162]<=8'd77;
		data_a[10163]<=8'd100;
		data_a[10164]<=8'd106;
		data_a[10165]<=8'd110;
		data_a[10166]<=8'd123;
		data_a[10167]<=8'd123;
		data_a[10168]<=8'd156;
		data_a[10169]<=8'd158;
		data_a[10170]<=8'd169;
		data_a[10171]<=8'd187;
		data_a[10172]<=8'd186;
		data_a[10173]<=8'd194;
		data_a[10174]<=8'd197;
		data_a[10175]<=8'd194;
		data_a[10176]<=8'd194;
		data_a[10177]<=8'd124;
		data_a[10178]<=8'd119;
		data_a[10179]<=8'd185;
		data_a[10180]<=8'd135;
		data_a[10181]<=8'd202;
		data_a[10182]<=8'd205;
		data_a[10183]<=8'd200;
		data_a[10184]<=8'd204;
		data_a[10185]<=8'd200;
		data_a[10186]<=8'd199;
		data_a[10187]<=8'd200;
		data_a[10188]<=8'd199;
		data_a[10189]<=8'd194;
		data_a[10190]<=8'd191;
		data_a[10191]<=8'd194;
		data_a[10192]<=8'd203;
		data_a[10193]<=8'd212;
		data_a[10194]<=8'd208;
		data_a[10195]<=8'd208;
		data_a[10196]<=8'd209;
		data_a[10197]<=8'd212;
		data_a[10198]<=8'd212;
		data_a[10199]<=8'd211;
		data_a[10200]<=8'd255;
		data_a[10201]<=8'd202;
		data_a[10202]<=8'd255;
		data_a[10203]<=8'd255;
		data_a[10204]<=8'd253;
		data_a[10205]<=8'd251;
		data_a[10206]<=8'd253;
		data_a[10207]<=8'd251;
		data_a[10208]<=8'd245;
		data_a[10209]<=8'd190;
		data_a[10210]<=8'd216;
		data_a[10211]<=8'd203;
		data_a[10212]<=8'd201;
		data_a[10213]<=8'd195;
		data_a[10214]<=8'd196;
		data_a[10215]<=8'd195;
		data_a[10216]<=8'd189;
		data_a[10217]<=8'd194;
		data_a[10218]<=8'd190;
		data_a[10219]<=8'd196;
		data_a[10220]<=8'd114;
		data_a[10221]<=8'd67;
		data_a[10222]<=8'd69;
		data_a[10223]<=8'd66;
		data_a[10224]<=8'd62;
		data_a[10225]<=8'd65;
		data_a[10226]<=8'd64;
		data_a[10227]<=8'd59;
		data_a[10228]<=8'd58;
		data_a[10229]<=8'd80;
		data_a[10230]<=8'd127;
		data_a[10231]<=8'd148;
		data_a[10232]<=8'd163;
		data_a[10233]<=8'd158;
		data_a[10234]<=8'd151;
		data_a[10235]<=8'd159;
		data_a[10236]<=8'd154;
		data_a[10237]<=8'd157;
		data_a[10238]<=8'd152;
		data_a[10239]<=8'd155;
		data_a[10240]<=8'd153;
		data_a[10241]<=8'd160;
		data_a[10242]<=8'd155;
		data_a[10243]<=8'd151;
		data_a[10244]<=8'd155;
		data_a[10245]<=8'd149;
		data_a[10246]<=8'd152;
		data_a[10247]<=8'd148;
		data_a[10248]<=8'd152;
		data_a[10249]<=8'd148;
		data_a[10250]<=8'd151;
		data_a[10251]<=8'd151;
		data_a[10252]<=8'd147;
		data_a[10253]<=8'd146;
		data_a[10254]<=8'd143;
		data_a[10255]<=8'd144;
		data_a[10256]<=8'd147;
		data_a[10257]<=8'd145;
		data_a[10258]<=8'd150;
		data_a[10259]<=8'd149;
		data_a[10260]<=8'd154;
		data_a[10261]<=8'd155;
		data_a[10262]<=8'd152;
		data_a[10263]<=8'd113;
		data_a[10264]<=8'd70;
		data_a[10265]<=8'd65;
		data_a[10266]<=8'd60;
		data_a[10267]<=8'd62;
		data_a[10268]<=8'd75;
		data_a[10269]<=8'd78;
		data_a[10270]<=8'd102;
		data_a[10271]<=8'd115;
		data_a[10272]<=8'd93;
		data_a[10273]<=8'd103;
		data_a[10274]<=8'd133;
		data_a[10275]<=8'd199;
		data_a[10276]<=8'd202;
		data_a[10277]<=8'd201;
		data_a[10278]<=8'd203;
		data_a[10279]<=8'd188;
		data_a[10280]<=8'd73;
		data_a[10281]<=8'd71;
		data_a[10282]<=8'd113;
		data_a[10283]<=8'd115;
		data_a[10284]<=8'd87;
		data_a[10285]<=8'd105;
		data_a[10286]<=8'd113;
		data_a[10287]<=8'd120;
		data_a[10288]<=8'd119;
		data_a[10289]<=8'd115;
		data_a[10290]<=8'd118;
		data_a[10291]<=8'd99;
		data_a[10292]<=8'd93;
		data_a[10293]<=8'd83;
		data_a[10294]<=8'd78;
		data_a[10295]<=8'd72;
		data_a[10296]<=8'd79;
		data_a[10297]<=8'd91;
		data_a[10298]<=8'd92;
		data_a[10299]<=8'd101;
		data_a[10300]<=8'd177;
		data_a[10301]<=8'd199;
		data_a[10302]<=8'd196;
		data_a[10303]<=8'd191;
		data_a[10304]<=8'd166;
		data_a[10305]<=8'd97;
		data_a[10306]<=8'd103;
		data_a[10307]<=8'd79;
		data_a[10308]<=8'd90;
		data_a[10309]<=8'd91;
		data_a[10310]<=8'd101;
		data_a[10311]<=8'd99;
		data_a[10312]<=8'd105;
		data_a[10313]<=8'd111;
		data_a[10314]<=8'd111;
		data_a[10315]<=8'd118;
		data_a[10316]<=8'd118;
		data_a[10317]<=8'd141;
		data_a[10318]<=8'd151;
		data_a[10319]<=8'd169;
		data_a[10320]<=8'd173;
		data_a[10321]<=8'd179;
		data_a[10322]<=8'd188;
		data_a[10323]<=8'd184;
		data_a[10324]<=8'd195;
		data_a[10325]<=8'd186;
		data_a[10326]<=8'd198;
		data_a[10327]<=8'd156;
		data_a[10328]<=8'd112;
		data_a[10329]<=8'd148;
		data_a[10330]<=8'd135;
		data_a[10331]<=8'd175;
		data_a[10332]<=8'd192;
		data_a[10333]<=8'd199;
		data_a[10334]<=8'd182;
		data_a[10335]<=8'd179;
		data_a[10336]<=8'd190;
		data_a[10337]<=8'd194;
		data_a[10338]<=8'd199;
		data_a[10339]<=8'd203;
		data_a[10340]<=8'd206;
		data_a[10341]<=8'd207;
		data_a[10342]<=8'd207;
		data_a[10343]<=8'd208;
		data_a[10344]<=8'd212;
		data_a[10345]<=8'd213;
		data_a[10346]<=8'd215;
		data_a[10347]<=8'd217;
		data_a[10348]<=8'd218;
		data_a[10349]<=8'd216;
		data_a[10350]<=8'd255;
		data_a[10351]<=8'd204;
		data_a[10352]<=8'd225;
		data_a[10353]<=8'd192;
		data_a[10354]<=8'd254;
		data_a[10355]<=8'd236;
		data_a[10356]<=8'd200;
		data_a[10357]<=8'd213;
		data_a[10358]<=8'd213;
		data_a[10359]<=8'd207;
		data_a[10360]<=8'd202;
		data_a[10361]<=8'd198;
		data_a[10362]<=8'd190;
		data_a[10363]<=8'd194;
		data_a[10364]<=8'd192;
		data_a[10365]<=8'd190;
		data_a[10366]<=8'd189;
		data_a[10367]<=8'd188;
		data_a[10368]<=8'd186;
		data_a[10369]<=8'd186;
		data_a[10370]<=8'd110;
		data_a[10371]<=8'd74;
		data_a[10372]<=8'd68;
		data_a[10373]<=8'd62;
		data_a[10374]<=8'd61;
		data_a[10375]<=8'd59;
		data_a[10376]<=8'd57;
		data_a[10377]<=8'd58;
		data_a[10378]<=8'd58;
		data_a[10379]<=8'd77;
		data_a[10380]<=8'd122;
		data_a[10381]<=8'd146;
		data_a[10382]<=8'd158;
		data_a[10383]<=8'd160;
		data_a[10384]<=8'd158;
		data_a[10385]<=8'd159;
		data_a[10386]<=8'd162;
		data_a[10387]<=8'd157;
		data_a[10388]<=8'd153;
		data_a[10389]<=8'd158;
		data_a[10390]<=8'd159;
		data_a[10391]<=8'd163;
		data_a[10392]<=8'd153;
		data_a[10393]<=8'd149;
		data_a[10394]<=8'd149;
		data_a[10395]<=8'd145;
		data_a[10396]<=8'd154;
		data_a[10397]<=8'd150;
		data_a[10398]<=8'd153;
		data_a[10399]<=8'd147;
		data_a[10400]<=8'd152;
		data_a[10401]<=8'd149;
		data_a[10402]<=8'd145;
		data_a[10403]<=8'd145;
		data_a[10404]<=8'd138;
		data_a[10405]<=8'd139;
		data_a[10406]<=8'd140;
		data_a[10407]<=8'd140;
		data_a[10408]<=8'd142;
		data_a[10409]<=8'd142;
		data_a[10410]<=8'd148;
		data_a[10411]<=8'd152;
		data_a[10412]<=8'd152;
		data_a[10413]<=8'd126;
		data_a[10414]<=8'd69;
		data_a[10415]<=8'd63;
		data_a[10416]<=8'd62;
		data_a[10417]<=8'd64;
		data_a[10418]<=8'd77;
		data_a[10419]<=8'd78;
		data_a[10420]<=8'd107;
		data_a[10421]<=8'd142;
		data_a[10422]<=8'd79;
		data_a[10423]<=8'd102;
		data_a[10424]<=8'd140;
		data_a[10425]<=8'd182;
		data_a[10426]<=8'd197;
		data_a[10427]<=8'd200;
		data_a[10428]<=8'd201;
		data_a[10429]<=8'd207;
		data_a[10430]<=8'd69;
		data_a[10431]<=8'd73;
		data_a[10432]<=8'd110;
		data_a[10433]<=8'd115;
		data_a[10434]<=8'd98;
		data_a[10435]<=8'd114;
		data_a[10436]<=8'd122;
		data_a[10437]<=8'd116;
		data_a[10438]<=8'd122;
		data_a[10439]<=8'd120;
		data_a[10440]<=8'd98;
		data_a[10441]<=8'd122;
		data_a[10442]<=8'd92;
		data_a[10443]<=8'd74;
		data_a[10444]<=8'd80;
		data_a[10445]<=8'd81;
		data_a[10446]<=8'd80;
		data_a[10447]<=8'd91;
		data_a[10448]<=8'd90;
		data_a[10449]<=8'd109;
		data_a[10450]<=8'd179;
		data_a[10451]<=8'd203;
		data_a[10452]<=8'd209;
		data_a[10453]<=8'd199;
		data_a[10454]<=8'd183;
		data_a[10455]<=8'd151;
		data_a[10456]<=8'd98;
		data_a[10457]<=8'd104;
		data_a[10458]<=8'd94;
		data_a[10459]<=8'd100;
		data_a[10460]<=8'd98;
		data_a[10461]<=8'd102;
		data_a[10462]<=8'd105;
		data_a[10463]<=8'd105;
		data_a[10464]<=8'd124;
		data_a[10465]<=8'd114;
		data_a[10466]<=8'd139;
		data_a[10467]<=8'd150;
		data_a[10468]<=8'd153;
		data_a[10469]<=8'd172;
		data_a[10470]<=8'd181;
		data_a[10471]<=8'd185;
		data_a[10472]<=8'd185;
		data_a[10473]<=8'd186;
		data_a[10474]<=8'd184;
		data_a[10475]<=8'd192;
		data_a[10476]<=8'd192;
		data_a[10477]<=8'd175;
		data_a[10478]<=8'd119;
		data_a[10479]<=8'd133;
		data_a[10480]<=8'd141;
		data_a[10481]<=8'd165;
		data_a[10482]<=8'd187;
		data_a[10483]<=8'd191;
		data_a[10484]<=8'd196;
		data_a[10485]<=8'd195;
		data_a[10486]<=8'd203;
		data_a[10487]<=8'd203;
		data_a[10488]<=8'd204;
		data_a[10489]<=8'd207;
		data_a[10490]<=8'd211;
		data_a[10491]<=8'd214;
		data_a[10492]<=8'd216;
		data_a[10493]<=8'd217;
		data_a[10494]<=8'd217;
		data_a[10495]<=8'd217;
		data_a[10496]<=8'd220;
		data_a[10497]<=8'd219;
		data_a[10498]<=8'd220;
		data_a[10499]<=8'd218;
		data_a[10500]<=8'd253;
		data_a[10501]<=8'd212;
		data_a[10502]<=8'd207;
		data_a[10503]<=8'd218;
		data_a[10504]<=8'd214;
		data_a[10505]<=8'd195;
		data_a[10506]<=8'd203;
		data_a[10507]<=8'd200;
		data_a[10508]<=8'd199;
		data_a[10509]<=8'd203;
		data_a[10510]<=8'd197;
		data_a[10511]<=8'd197;
		data_a[10512]<=8'd195;
		data_a[10513]<=8'd193;
		data_a[10514]<=8'd194;
		data_a[10515]<=8'd189;
		data_a[10516]<=8'd185;
		data_a[10517]<=8'd186;
		data_a[10518]<=8'd186;
		data_a[10519]<=8'd174;
		data_a[10520]<=8'd86;
		data_a[10521]<=8'd84;
		data_a[10522]<=8'd61;
		data_a[10523]<=8'd64;
		data_a[10524]<=8'd63;
		data_a[10525]<=8'd61;
		data_a[10526]<=8'd60;
		data_a[10527]<=8'd65;
		data_a[10528]<=8'd64;
		data_a[10529]<=8'd81;
		data_a[10530]<=8'd123;
		data_a[10531]<=8'd148;
		data_a[10532]<=8'd155;
		data_a[10533]<=8'd162;
		data_a[10534]<=8'd162;
		data_a[10535]<=8'd161;
		data_a[10536]<=8'd165;
		data_a[10537]<=8'd159;
		data_a[10538]<=8'd156;
		data_a[10539]<=8'd162;
		data_a[10540]<=8'd161;
		data_a[10541]<=8'd158;
		data_a[10542]<=8'd151;
		data_a[10543]<=8'd144;
		data_a[10544]<=8'd143;
		data_a[10545]<=8'd143;
		data_a[10546]<=8'd154;
		data_a[10547]<=8'd154;
		data_a[10548]<=8'd155;
		data_a[10549]<=8'd151;
		data_a[10550]<=8'd152;
		data_a[10551]<=8'd150;
		data_a[10552]<=8'd148;
		data_a[10553]<=8'd146;
		data_a[10554]<=8'd142;
		data_a[10555]<=8'd138;
		data_a[10556]<=8'd136;
		data_a[10557]<=8'd138;
		data_a[10558]<=8'd142;
		data_a[10559]<=8'd149;
		data_a[10560]<=8'd155;
		data_a[10561]<=8'd152;
		data_a[10562]<=8'd145;
		data_a[10563]<=8'd134;
		data_a[10564]<=8'd72;
		data_a[10565]<=8'd72;
		data_a[10566]<=8'd59;
		data_a[10567]<=8'd62;
		data_a[10568]<=8'd68;
		data_a[10569]<=8'd64;
		data_a[10570]<=8'd137;
		data_a[10571]<=8'd126;
		data_a[10572]<=8'd77;
		data_a[10573]<=8'd90;
		data_a[10574]<=8'd110;
		data_a[10575]<=8'd193;
		data_a[10576]<=8'd200;
		data_a[10577]<=8'd196;
		data_a[10578]<=8'd199;
		data_a[10579]<=8'd204;
		data_a[10580]<=8'd70;
		data_a[10581]<=8'd70;
		data_a[10582]<=8'd110;
		data_a[10583]<=8'd116;
		data_a[10584]<=8'd100;
		data_a[10585]<=8'd117;
		data_a[10586]<=8'd122;
		data_a[10587]<=8'd114;
		data_a[10588]<=8'd113;
		data_a[10589]<=8'd111;
		data_a[10590]<=8'd113;
		data_a[10591]<=8'd73;
		data_a[10592]<=8'd66;
		data_a[10593]<=8'd65;
		data_a[10594]<=8'd68;
		data_a[10595]<=8'd81;
		data_a[10596]<=8'd85;
		data_a[10597]<=8'd88;
		data_a[10598]<=8'd89;
		data_a[10599]<=8'd126;
		data_a[10600]<=8'd174;
		data_a[10601]<=8'd208;
		data_a[10602]<=8'd222;
		data_a[10603]<=8'd199;
		data_a[10604]<=8'd200;
		data_a[10605]<=8'd168;
		data_a[10606]<=8'd119;
		data_a[10607]<=8'd99;
		data_a[10608]<=8'd99;
		data_a[10609]<=8'd92;
		data_a[10610]<=8'd91;
		data_a[10611]<=8'd110;
		data_a[10612]<=8'd111;
		data_a[10613]<=8'd102;
		data_a[10614]<=8'd124;
		data_a[10615]<=8'd130;
		data_a[10616]<=8'd133;
		data_a[10617]<=8'd155;
		data_a[10618]<=8'd171;
		data_a[10619]<=8'd184;
		data_a[10620]<=8'd188;
		data_a[10621]<=8'd188;
		data_a[10622]<=8'd189;
		data_a[10623]<=8'd184;
		data_a[10624]<=8'd187;
		data_a[10625]<=8'd186;
		data_a[10626]<=8'd190;
		data_a[10627]<=8'd173;
		data_a[10628]<=8'd116;
		data_a[10629]<=8'd146;
		data_a[10630]<=8'd136;
		data_a[10631]<=8'd149;
		data_a[10632]<=8'd202;
		data_a[10633]<=8'd204;
		data_a[10634]<=8'd198;
		data_a[10635]<=8'd204;
		data_a[10636]<=8'd204;
		data_a[10637]<=8'd207;
		data_a[10638]<=8'd210;
		data_a[10639]<=8'd211;
		data_a[10640]<=8'd212;
		data_a[10641]<=8'd212;
		data_a[10642]<=8'd214;
		data_a[10643]<=8'd215;
		data_a[10644]<=8'd217;
		data_a[10645]<=8'd217;
		data_a[10646]<=8'd220;
		data_a[10647]<=8'd219;
		data_a[10648]<=8'd223;
		data_a[10649]<=8'd222;
		data_a[10650]<=8'd253;
		data_a[10651]<=8'd205;
		data_a[10652]<=8'd204;
		data_a[10653]<=8'd205;
		data_a[10654]<=8'd207;
		data_a[10655]<=8'd207;
		data_a[10656]<=8'd205;
		data_a[10657]<=8'd178;
		data_a[10658]<=8'd198;
		data_a[10659]<=8'd202;
		data_a[10660]<=8'd199;
		data_a[10661]<=8'd192;
		data_a[10662]<=8'd191;
		data_a[10663]<=8'd190;
		data_a[10664]<=8'd186;
		data_a[10665]<=8'd189;
		data_a[10666]<=8'd186;
		data_a[10667]<=8'd182;
		data_a[10668]<=8'd182;
		data_a[10669]<=8'd156;
		data_a[10670]<=8'd82;
		data_a[10671]<=8'd68;
		data_a[10672]<=8'd62;
		data_a[10673]<=8'd60;
		data_a[10674]<=8'd58;
		data_a[10675]<=8'd60;
		data_a[10676]<=8'd60;
		data_a[10677]<=8'd65;
		data_a[10678]<=8'd64;
		data_a[10679]<=8'd83;
		data_a[10680]<=8'd123;
		data_a[10681]<=8'd143;
		data_a[10682]<=8'd156;
		data_a[10683]<=8'd160;
		data_a[10684]<=8'd158;
		data_a[10685]<=8'd164;
		data_a[10686]<=8'd159;
		data_a[10687]<=8'd165;
		data_a[10688]<=8'd162;
		data_a[10689]<=8'd165;
		data_a[10690]<=8'd163;
		data_a[10691]<=8'd157;
		data_a[10692]<=8'd159;
		data_a[10693]<=8'd153;
		data_a[10694]<=8'd152;
		data_a[10695]<=8'd154;
		data_a[10696]<=8'd160;
		data_a[10697]<=8'd161;
		data_a[10698]<=8'd156;
		data_a[10699]<=8'd155;
		data_a[10700]<=8'd150;
		data_a[10701]<=8'd152;
		data_a[10702]<=8'd149;
		data_a[10703]<=8'd146;
		data_a[10704]<=8'd147;
		data_a[10705]<=8'd139;
		data_a[10706]<=8'd137;
		data_a[10707]<=8'd143;
		data_a[10708]<=8'd144;
		data_a[10709]<=8'd146;
		data_a[10710]<=8'd151;
		data_a[10711]<=8'd150;
		data_a[10712]<=8'd142;
		data_a[10713]<=8'd138;
		data_a[10714]<=8'd83;
		data_a[10715]<=8'd61;
		data_a[10716]<=8'd67;
		data_a[10717]<=8'd63;
		data_a[10718]<=8'd68;
		data_a[10719]<=8'd76;
		data_a[10720]<=8'd80;
		data_a[10721]<=8'd98;
		data_a[10722]<=8'd76;
		data_a[10723]<=8'd85;
		data_a[10724]<=8'd109;
		data_a[10725]<=8'd191;
		data_a[10726]<=8'd200;
		data_a[10727]<=8'd198;
		data_a[10728]<=8'd202;
		data_a[10729]<=8'd203;
		data_a[10730]<=8'd78;
		data_a[10731]<=8'd69;
		data_a[10732]<=8'd121;
		data_a[10733]<=8'd123;
		data_a[10734]<=8'd102;
		data_a[10735]<=8'd120;
		data_a[10736]<=8'd115;
		data_a[10737]<=8'd111;
		data_a[10738]<=8'd102;
		data_a[10739]<=8'd124;
		data_a[10740]<=8'd62;
		data_a[10741]<=8'd70;
		data_a[10742]<=8'd71;
		data_a[10743]<=8'd76;
		data_a[10744]<=8'd72;
		data_a[10745]<=8'd90;
		data_a[10746]<=8'd67;
		data_a[10747]<=8'd90;
		data_a[10748]<=8'd98;
		data_a[10749]<=8'd144;
		data_a[10750]<=8'd172;
		data_a[10751]<=8'd202;
		data_a[10752]<=8'd221;
		data_a[10753]<=8'd207;
		data_a[10754]<=8'd205;
		data_a[10755]<=8'd175;
		data_a[10756]<=8'd155;
		data_a[10757]<=8'd107;
		data_a[10758]<=8'd101;
		data_a[10759]<=8'd102;
		data_a[10760]<=8'd107;
		data_a[10761]<=8'd104;
		data_a[10762]<=8'd113;
		data_a[10763]<=8'd115;
		data_a[10764]<=8'd124;
		data_a[10765]<=8'd124;
		data_a[10766]<=8'd143;
		data_a[10767]<=8'd165;
		data_a[10768]<=8'd173;
		data_a[10769]<=8'd185;
		data_a[10770]<=8'd186;
		data_a[10771]<=8'd187;
		data_a[10772]<=8'd182;
		data_a[10773]<=8'd186;
		data_a[10774]<=8'd184;
		data_a[10775]<=8'd182;
		data_a[10776]<=8'd191;
		data_a[10777]<=8'd173;
		data_a[10778]<=8'd113;
		data_a[10779]<=8'd136;
		data_a[10780]<=8'd193;
		data_a[10781]<=8'd148;
		data_a[10782]<=8'd216;
		data_a[10783]<=8'd200;
		data_a[10784]<=8'd209;
		data_a[10785]<=8'd205;
		data_a[10786]<=8'd208;
		data_a[10787]<=8'd209;
		data_a[10788]<=8'd210;
		data_a[10789]<=8'd211;
		data_a[10790]<=8'd214;
		data_a[10791]<=8'd216;
		data_a[10792]<=8'd219;
		data_a[10793]<=8'd221;
		data_a[10794]<=8'd221;
		data_a[10795]<=8'd219;
		data_a[10796]<=8'd221;
		data_a[10797]<=8'd219;
		data_a[10798]<=8'd225;
		data_a[10799]<=8'd224;
		data_a[10800]<=8'd255;
		data_a[10801]<=8'd196;
		data_a[10802]<=8'd201;
		data_a[10803]<=8'd204;
		data_a[10804]<=8'd204;
		data_a[10805]<=8'd199;
		data_a[10806]<=8'd200;
		data_a[10807]<=8'd200;
		data_a[10808]<=8'd192;
		data_a[10809]<=8'd183;
		data_a[10810]<=8'd197;
		data_a[10811]<=8'd192;
		data_a[10812]<=8'd186;
		data_a[10813]<=8'd187;
		data_a[10814]<=8'd187;
		data_a[10815]<=8'd185;
		data_a[10816]<=8'd183;
		data_a[10817]<=8'd181;
		data_a[10818]<=8'd174;
		data_a[10819]<=8'd121;
		data_a[10820]<=8'd74;
		data_a[10821]<=8'd67;
		data_a[10822]<=8'd67;
		data_a[10823]<=8'd67;
		data_a[10824]<=8'd63;
		data_a[10825]<=8'd63;
		data_a[10826]<=8'd56;
		data_a[10827]<=8'd60;
		data_a[10828]<=8'd66;
		data_a[10829]<=8'd80;
		data_a[10830]<=8'd115;
		data_a[10831]<=8'd153;
		data_a[10832]<=8'd157;
		data_a[10833]<=8'd161;
		data_a[10834]<=8'd168;
		data_a[10835]<=8'd163;
		data_a[10836]<=8'd163;
		data_a[10837]<=8'd165;
		data_a[10838]<=8'd167;
		data_a[10839]<=8'd165;
		data_a[10840]<=8'd171;
		data_a[10841]<=8'd158;
		data_a[10842]<=8'd167;
		data_a[10843]<=8'd159;
		data_a[10844]<=8'd165;
		data_a[10845]<=8'd159;
		data_a[10846]<=8'd164;
		data_a[10847]<=8'd164;
		data_a[10848]<=8'd155;
		data_a[10849]<=8'd156;
		data_a[10850]<=8'd160;
		data_a[10851]<=8'd152;
		data_a[10852]<=8'd157;
		data_a[10853]<=8'd102;
		data_a[10854]<=8'd143;
		data_a[10855]<=8'd145;
		data_a[10856]<=8'd141;
		data_a[10857]<=8'd140;
		data_a[10858]<=8'd144;
		data_a[10859]<=8'd149;
		data_a[10860]<=8'd152;
		data_a[10861]<=8'd151;
		data_a[10862]<=8'd143;
		data_a[10863]<=8'd132;
		data_a[10864]<=8'd85;
		data_a[10865]<=8'd61;
		data_a[10866]<=8'd62;
		data_a[10867]<=8'd65;
		data_a[10868]<=8'd65;
		data_a[10869]<=8'd67;
		data_a[10870]<=8'd80;
		data_a[10871]<=8'd92;
		data_a[10872]<=8'd74;
		data_a[10873]<=8'd95;
		data_a[10874]<=8'd121;
		data_a[10875]<=8'd188;
		data_a[10876]<=8'd198;
		data_a[10877]<=8'd199;
		data_a[10878]<=8'd200;
		data_a[10879]<=8'd195;
		data_a[10880]<=8'd58;
		data_a[10881]<=8'd73;
		data_a[10882]<=8'd111;
		data_a[10883]<=8'd108;
		data_a[10884]<=8'd113;
		data_a[10885]<=8'd118;
		data_a[10886]<=8'd110;
		data_a[10887]<=8'd107;
		data_a[10888]<=8'd119;
		data_a[10889]<=8'd70;
		data_a[10890]<=8'd85;
		data_a[10891]<=8'd72;
		data_a[10892]<=8'd76;
		data_a[10893]<=8'd74;
		data_a[10894]<=8'd69;
		data_a[10895]<=8'd101;
		data_a[10896]<=8'd81;
		data_a[10897]<=8'd85;
		data_a[10898]<=8'd90;
		data_a[10899]<=8'd150;
		data_a[10900]<=8'd173;
		data_a[10901]<=8'd203;
		data_a[10902]<=8'd208;
		data_a[10903]<=8'd213;
		data_a[10904]<=8'd205;
		data_a[10905]<=8'd182;
		data_a[10906]<=8'd163;
		data_a[10907]<=8'd135;
		data_a[10908]<=8'd111;
		data_a[10909]<=8'd105;
		data_a[10910]<=8'd109;
		data_a[10911]<=8'd115;
		data_a[10912]<=8'd116;
		data_a[10913]<=8'd124;
		data_a[10914]<=8'd132;
		data_a[10915]<=8'd146;
		data_a[10916]<=8'd164;
		data_a[10917]<=8'd175;
		data_a[10918]<=8'd181;
		data_a[10919]<=8'd188;
		data_a[10920]<=8'd187;
		data_a[10921]<=8'd185;
		data_a[10922]<=8'd185;
		data_a[10923]<=8'd186;
		data_a[10924]<=8'd181;
		data_a[10925]<=8'd177;
		data_a[10926]<=8'd185;
		data_a[10927]<=8'd171;
		data_a[10928]<=8'd126;
		data_a[10929]<=8'd130;
		data_a[10930]<=8'd227;
		data_a[10931]<=8'd130;
		data_a[10932]<=8'd220;
		data_a[10933]<=8'd206;
		data_a[10934]<=8'd210;
		data_a[10935]<=8'd209;
		data_a[10936]<=8'd212;
		data_a[10937]<=8'd213;
		data_a[10938]<=8'd213;
		data_a[10939]<=8'd214;
		data_a[10940]<=8'd215;
		data_a[10941]<=8'd217;
		data_a[10942]<=8'd219;
		data_a[10943]<=8'd220;
		data_a[10944]<=8'd222;
		data_a[10945]<=8'd222;
		data_a[10946]<=8'd223;
		data_a[10947]<=8'd224;
		data_a[10948]<=8'd225;
		data_a[10949]<=8'd225;
		data_a[10950]<=8'd255;
		data_a[10951]<=8'd194;
		data_a[10952]<=8'd195;
		data_a[10953]<=8'd193;
		data_a[10954]<=8'd196;
		data_a[10955]<=8'd198;
		data_a[10956]<=8'd196;
		data_a[10957]<=8'd188;
		data_a[10958]<=8'd181;
		data_a[10959]<=8'd198;
		data_a[10960]<=8'd176;
		data_a[10961]<=8'd182;
		data_a[10962]<=8'd180;
		data_a[10963]<=8'd181;
		data_a[10964]<=8'd184;
		data_a[10965]<=8'd185;
		data_a[10966]<=8'd182;
		data_a[10967]<=8'd185;
		data_a[10968]<=8'd169;
		data_a[10969]<=8'd85;
		data_a[10970]<=8'd67;
		data_a[10971]<=8'd70;
		data_a[10972]<=8'd65;
		data_a[10973]<=8'd62;
		data_a[10974]<=8'd64;
		data_a[10975]<=8'd57;
		data_a[10976]<=8'd53;
		data_a[10977]<=8'd58;
		data_a[10978]<=8'd65;
		data_a[10979]<=8'd81;
		data_a[10980]<=8'd117;
		data_a[10981]<=8'd145;
		data_a[10982]<=8'd161;
		data_a[10983]<=8'd160;
		data_a[10984]<=8'd159;
		data_a[10985]<=8'd170;
		data_a[10986]<=8'd167;
		data_a[10987]<=8'd163;
		data_a[10988]<=8'd168;
		data_a[10989]<=8'd174;
		data_a[10990]<=8'd157;
		data_a[10991]<=8'd163;
		data_a[10992]<=8'd168;
		data_a[10993]<=8'd166;
		data_a[10994]<=8'd172;
		data_a[10995]<=8'd159;
		data_a[10996]<=8'd157;
		data_a[10997]<=8'd160;
		data_a[10998]<=8'd160;
		data_a[10999]<=8'd166;
		data_a[11000]<=8'd151;
		data_a[11001]<=8'd164;
		data_a[11002]<=8'd158;
		data_a[11003]<=8'd152;
		data_a[11004]<=8'd156;
		data_a[11005]<=8'd152;
		data_a[11006]<=8'd146;
		data_a[11007]<=8'd145;
		data_a[11008]<=8'd147;
		data_a[11009]<=8'd150;
		data_a[11010]<=8'd151;
		data_a[11011]<=8'd150;
		data_a[11012]<=8'd143;
		data_a[11013]<=8'd133;
		data_a[11014]<=8'd92;
		data_a[11015]<=8'd63;
		data_a[11016]<=8'd64;
		data_a[11017]<=8'd65;
		data_a[11018]<=8'd69;
		data_a[11019]<=8'd71;
		data_a[11020]<=8'd72;
		data_a[11021]<=8'd77;
		data_a[11022]<=8'd93;
		data_a[11023]<=8'd91;
		data_a[11024]<=8'd158;
		data_a[11025]<=8'd189;
		data_a[11026]<=8'd197;
		data_a[11027]<=8'd197;
		data_a[11028]<=8'd191;
		data_a[11029]<=8'd188;
		data_a[11030]<=8'd68;
		data_a[11031]<=8'd71;
		data_a[11032]<=8'd118;
		data_a[11033]<=8'd126;
		data_a[11034]<=8'd126;
		data_a[11035]<=8'd115;
		data_a[11036]<=8'd109;
		data_a[11037]<=8'd94;
		data_a[11038]<=8'd85;
		data_a[11039]<=8'd71;
		data_a[11040]<=8'd102;
		data_a[11041]<=8'd60;
		data_a[11042]<=8'd86;
		data_a[11043]<=8'd76;
		data_a[11044]<=8'd71;
		data_a[11045]<=8'd88;
		data_a[11046]<=8'd87;
		data_a[11047]<=8'd104;
		data_a[11048]<=8'd101;
		data_a[11049]<=8'd150;
		data_a[11050]<=8'd164;
		data_a[11051]<=8'd201;
		data_a[11052]<=8'd210;
		data_a[11053]<=8'd215;
		data_a[11054]<=8'd208;
		data_a[11055]<=8'd185;
		data_a[11056]<=8'd170;
		data_a[11057]<=8'd148;
		data_a[11058]<=8'd124;
		data_a[11059]<=8'd128;
		data_a[11060]<=8'd132;
		data_a[11061]<=8'd127;
		data_a[11062]<=8'd134;
		data_a[11063]<=8'd141;
		data_a[11064]<=8'd151;
		data_a[11065]<=8'd159;
		data_a[11066]<=8'd167;
		data_a[11067]<=8'd174;
		data_a[11068]<=8'd184;
		data_a[11069]<=8'd193;
		data_a[11070]<=8'd182;
		data_a[11071]<=8'd187;
		data_a[11072]<=8'd183;
		data_a[11073]<=8'd174;
		data_a[11074]<=8'd183;
		data_a[11075]<=8'd178;
		data_a[11076]<=8'd184;
		data_a[11077]<=8'd174;
		data_a[11078]<=8'd117;
		data_a[11079]<=8'd119;
		data_a[11080]<=8'd186;
		data_a[11081]<=8'd189;
		data_a[11082]<=8'd194;
		data_a[11083]<=8'd211;
		data_a[11084]<=8'd214;
		data_a[11085]<=8'd213;
		data_a[11086]<=8'd214;
		data_a[11087]<=8'd215;
		data_a[11088]<=8'd217;
		data_a[11089]<=8'd219;
		data_a[11090]<=8'd220;
		data_a[11091]<=8'd221;
		data_a[11092]<=8'd222;
		data_a[11093]<=8'd222;
		data_a[11094]<=8'd224;
		data_a[11095]<=8'd225;
		data_a[11096]<=8'd226;
		data_a[11097]<=8'd227;
		data_a[11098]<=8'd229;
		data_a[11099]<=8'd229;
		data_a[11100]<=8'd251;
		data_a[11101]<=8'd188;
		data_a[11102]<=8'd194;
		data_a[11103]<=8'd193;
		data_a[11104]<=8'd187;
		data_a[11105]<=8'd181;
		data_a[11106]<=8'd186;
		data_a[11107]<=8'd192;
		data_a[11108]<=8'd187;
		data_a[11109]<=8'd182;
		data_a[11110]<=8'd181;
		data_a[11111]<=8'd190;
		data_a[11112]<=8'd161;
		data_a[11113]<=8'd179;
		data_a[11114]<=8'd184;
		data_a[11115]<=8'd183;
		data_a[11116]<=8'd178;
		data_a[11117]<=8'd185;
		data_a[11118]<=8'd90;
		data_a[11119]<=8'd100;
		data_a[11120]<=8'd65;
		data_a[11121]<=8'd66;
		data_a[11122]<=8'd67;
		data_a[11123]<=8'd66;
		data_a[11124]<=8'd63;
		data_a[11125]<=8'd51;
		data_a[11126]<=8'd54;
		data_a[11127]<=8'd58;
		data_a[11128]<=8'd65;
		data_a[11129]<=8'd79;
		data_a[11130]<=8'd120;
		data_a[11131]<=8'd142;
		data_a[11132]<=8'd162;
		data_a[11133]<=8'd170;
		data_a[11134]<=8'd171;
		data_a[11135]<=8'd169;
		data_a[11136]<=8'd173;
		data_a[11137]<=8'd173;
		data_a[11138]<=8'd168;
		data_a[11139]<=8'd172;
		data_a[11140]<=8'd170;
		data_a[11141]<=8'd172;
		data_a[11142]<=8'd170;
		data_a[11143]<=8'd172;
		data_a[11144]<=8'd167;
		data_a[11145]<=8'd157;
		data_a[11146]<=8'd162;
		data_a[11147]<=8'd161;
		data_a[11148]<=8'd155;
		data_a[11149]<=8'd163;
		data_a[11150]<=8'd171;
		data_a[11151]<=8'd166;
		data_a[11152]<=8'd169;
		data_a[11153]<=8'd163;
		data_a[11154]<=8'd165;
		data_a[11155]<=8'd158;
		data_a[11156]<=8'd153;
		data_a[11157]<=8'd151;
		data_a[11158]<=8'd150;
		data_a[11159]<=8'd150;
		data_a[11160]<=8'd150;
		data_a[11161]<=8'd151;
		data_a[11162]<=8'd144;
		data_a[11163]<=8'd134;
		data_a[11164]<=8'd88;
		data_a[11165]<=8'd62;
		data_a[11166]<=8'd63;
		data_a[11167]<=8'd63;
		data_a[11168]<=8'd68;
		data_a[11169]<=8'd74;
		data_a[11170]<=8'd77;
		data_a[11171]<=8'd85;
		data_a[11172]<=8'd91;
		data_a[11173]<=8'd101;
		data_a[11174]<=8'd153;
		data_a[11175]<=8'd184;
		data_a[11176]<=8'd189;
		data_a[11177]<=8'd201;
		data_a[11178]<=8'd201;
		data_a[11179]<=8'd193;
		data_a[11180]<=8'd89;
		data_a[11181]<=8'd67;
		data_a[11182]<=8'd136;
		data_a[11183]<=8'd133;
		data_a[11184]<=8'd126;
		data_a[11185]<=8'd123;
		data_a[11186]<=8'd115;
		data_a[11187]<=8'd89;
		data_a[11188]<=8'd62;
		data_a[11189]<=8'd110;
		data_a[11190]<=8'd115;
		data_a[11191]<=8'd96;
		data_a[11192]<=8'd91;
		data_a[11193]<=8'd65;
		data_a[11194]<=8'd71;
		data_a[11195]<=8'd94;
		data_a[11196]<=8'd99;
		data_a[11197]<=8'd101;
		data_a[11198]<=8'd108;
		data_a[11199]<=8'd158;
		data_a[11200]<=8'd161;
		data_a[11201]<=8'd188;
		data_a[11202]<=8'd208;
		data_a[11203]<=8'd214;
		data_a[11204]<=8'd214;
		data_a[11205]<=8'd214;
		data_a[11206]<=8'd179;
		data_a[11207]<=8'd162;
		data_a[11208]<=8'd148;
		data_a[11209]<=8'd141;
		data_a[11210]<=8'd147;
		data_a[11211]<=8'd151;
		data_a[11212]<=8'd158;
		data_a[11213]<=8'd160;
		data_a[11214]<=8'd168;
		data_a[11215]<=8'd176;
		data_a[11216]<=8'd181;
		data_a[11217]<=8'd188;
		data_a[11218]<=8'd197;
		data_a[11219]<=8'd202;
		data_a[11220]<=8'd193;
		data_a[11221]<=8'd187;
		data_a[11222]<=8'd179;
		data_a[11223]<=8'd185;
		data_a[11224]<=8'd178;
		data_a[11225]<=8'd177;
		data_a[11226]<=8'd180;
		data_a[11227]<=8'd174;
		data_a[11228]<=8'd118;
		data_a[11229]<=8'd117;
		data_a[11230]<=8'd149;
		data_a[11231]<=8'd208;
		data_a[11232]<=8'd182;
		data_a[11233]<=8'd211;
		data_a[11234]<=8'd214;
		data_a[11235]<=8'd216;
		data_a[11236]<=8'd216;
		data_a[11237]<=8'd217;
		data_a[11238]<=8'd219;
		data_a[11239]<=8'd221;
		data_a[11240]<=8'd222;
		data_a[11241]<=8'd223;
		data_a[11242]<=8'd224;
		data_a[11243]<=8'd225;
		data_a[11244]<=8'd224;
		data_a[11245]<=8'd225;
		data_a[11246]<=8'd226;
		data_a[11247]<=8'd227;
		data_a[11248]<=8'd227;
		data_a[11249]<=8'd228;
		data_a[11250]<=8'd255;
		data_a[11251]<=8'd178;
		data_a[11252]<=8'd176;
		data_a[11253]<=8'd184;
		data_a[11254]<=8'd191;
		data_a[11255]<=8'd189;
		data_a[11256]<=8'd185;
		data_a[11257]<=8'd184;
		data_a[11258]<=8'd188;
		data_a[11259]<=8'd179;
		data_a[11260]<=8'd184;
		data_a[11261]<=8'd180;
		data_a[11262]<=8'd182;
		data_a[11263]<=8'd184;
		data_a[11264]<=8'd150;
		data_a[11265]<=8'd164;
		data_a[11266]<=8'd148;
		data_a[11267]<=8'd179;
		data_a[11268]<=8'd84;
		data_a[11269]<=8'd102;
		data_a[11270]<=8'd68;
		data_a[11271]<=8'd66;
		data_a[11272]<=8'd72;
		data_a[11273]<=8'd66;
		data_a[11274]<=8'd55;
		data_a[11275]<=8'd50;
		data_a[11276]<=8'd58;
		data_a[11277]<=8'd57;
		data_a[11278]<=8'd64;
		data_a[11279]<=8'd75;
		data_a[11280]<=8'd123;
		data_a[11281]<=8'd148;
		data_a[11282]<=8'd160;
		data_a[11283]<=8'd161;
		data_a[11284]<=8'd172;
		data_a[11285]<=8'd176;
		data_a[11286]<=8'd181;
		data_a[11287]<=8'd179;
		data_a[11288]<=8'd172;
		data_a[11289]<=8'd170;
		data_a[11290]<=8'd168;
		data_a[11291]<=8'd162;
		data_a[11292]<=8'd161;
		data_a[11293]<=8'd163;
		data_a[11294]<=8'd160;
		data_a[11295]<=8'd157;
		data_a[11296]<=8'd162;
		data_a[11297]<=8'd157;
		data_a[11298]<=8'd165;
		data_a[11299]<=8'd163;
		data_a[11300]<=8'd166;
		data_a[11301]<=8'd160;
		data_a[11302]<=8'd163;
		data_a[11303]<=8'd161;
		data_a[11304]<=8'd166;
		data_a[11305]<=8'd168;
		data_a[11306]<=8'd157;
		data_a[11307]<=8'd154;
		data_a[11308]<=8'd150;
		data_a[11309]<=8'd147;
		data_a[11310]<=8'd147;
		data_a[11311]<=8'd150;
		data_a[11312]<=8'd144;
		data_a[11313]<=8'd133;
		data_a[11314]<=8'd92;
		data_a[11315]<=8'd70;
		data_a[11316]<=8'd65;
		data_a[11317]<=8'd62;
		data_a[11318]<=8'd64;
		data_a[11319]<=8'd68;
		data_a[11320]<=8'd77;
		data_a[11321]<=8'd85;
		data_a[11322]<=8'd90;
		data_a[11323]<=8'd125;
		data_a[11324]<=8'd178;
		data_a[11325]<=8'd185;
		data_a[11326]<=8'd199;
		data_a[11327]<=8'd199;
		data_a[11328]<=8'd191;
		data_a[11329]<=8'd200;
		data_a[11330]<=8'd162;
		data_a[11331]<=8'd77;
		data_a[11332]<=8'd125;
		data_a[11333]<=8'd133;
		data_a[11334]<=8'd129;
		data_a[11335]<=8'd113;
		data_a[11336]<=8'd108;
		data_a[11337]<=8'd77;
		data_a[11338]<=8'd69;
		data_a[11339]<=8'd102;
		data_a[11340]<=8'd134;
		data_a[11341]<=8'd67;
		data_a[11342]<=8'd85;
		data_a[11343]<=8'd91;
		data_a[11344]<=8'd85;
		data_a[11345]<=8'd99;
		data_a[11346]<=8'd100;
		data_a[11347]<=8'd107;
		data_a[11348]<=8'd121;
		data_a[11349]<=8'd147;
		data_a[11350]<=8'd166;
		data_a[11351]<=8'd189;
		data_a[11352]<=8'd209;
		data_a[11353]<=8'd218;
		data_a[11354]<=8'd210;
		data_a[11355]<=8'd226;
		data_a[11356]<=8'd185;
		data_a[11357]<=8'd171;
		data_a[11358]<=8'd154;
		data_a[11359]<=8'd146;
		data_a[11360]<=8'd159;
		data_a[11361]<=8'd156;
		data_a[11362]<=8'd163;
		data_a[11363]<=8'd163;
		data_a[11364]<=8'd171;
		data_a[11365]<=8'd180;
		data_a[11366]<=8'd185;
		data_a[11367]<=8'd192;
		data_a[11368]<=8'd199;
		data_a[11369]<=8'd201;
		data_a[11370]<=8'd203;
		data_a[11371]<=8'd188;
		data_a[11372]<=8'd189;
		data_a[11373]<=8'd187;
		data_a[11374]<=8'd184;
		data_a[11375]<=8'd172;
		data_a[11376]<=8'd180;
		data_a[11377]<=8'd169;
		data_a[11378]<=8'd125;
		data_a[11379]<=8'd111;
		data_a[11380]<=8'd122;
		data_a[11381]<=8'd182;
		data_a[11382]<=8'd165;
		data_a[11383]<=8'd212;
		data_a[11384]<=8'd218;
		data_a[11385]<=8'd216;
		data_a[11386]<=8'd219;
		data_a[11387]<=8'd219;
		data_a[11388]<=8'd219;
		data_a[11389]<=8'd221;
		data_a[11390]<=8'd222;
		data_a[11391]<=8'd223;
		data_a[11392]<=8'd225;
		data_a[11393]<=8'd227;
		data_a[11394]<=8'd227;
		data_a[11395]<=8'd227;
		data_a[11396]<=8'd228;
		data_a[11397]<=8'd229;
		data_a[11398]<=8'd229;
		data_a[11399]<=8'd229;
		data_a[11400]<=8'd254;
		data_a[11401]<=8'd178;
		data_a[11402]<=8'd181;
		data_a[11403]<=8'd182;
		data_a[11404]<=8'd183;
		data_a[11405]<=8'd186;
		data_a[11406]<=8'd185;
		data_a[11407]<=8'd183;
		data_a[11408]<=8'd185;
		data_a[11409]<=8'd177;
		data_a[11410]<=8'd183;
		data_a[11411]<=8'd182;
		data_a[11412]<=8'd177;
		data_a[11413]<=8'd176;
		data_a[11414]<=8'd176;
		data_a[11415]<=8'd185;
		data_a[11416]<=8'd152;
		data_a[11417]<=8'd164;
		data_a[11418]<=8'd94;
		data_a[11419]<=8'd85;
		data_a[11420]<=8'd99;
		data_a[11421]<=8'd68;
		data_a[11422]<=8'd67;
		data_a[11423]<=8'd69;
		data_a[11424]<=8'd49;
		data_a[11425]<=8'd50;
		data_a[11426]<=8'd59;
		data_a[11427]<=8'd53;
		data_a[11428]<=8'd63;
		data_a[11429]<=8'd75;
		data_a[11430]<=8'd124;
		data_a[11431]<=8'd155;
		data_a[11432]<=8'd161;
		data_a[11433]<=8'd174;
		data_a[11434]<=8'd173;
		data_a[11435]<=8'd192;
		data_a[11436]<=8'd169;
		data_a[11437]<=8'd172;
		data_a[11438]<=8'd169;
		data_a[11439]<=8'd151;
		data_a[11440]<=8'd152;
		data_a[11441]<=8'd150;
		data_a[11442]<=8'd149;
		data_a[11443]<=8'd142;
		data_a[11444]<=8'd152;
		data_a[11445]<=8'd150;
		data_a[11446]<=8'd148;
		data_a[11447]<=8'd151;
		data_a[11448]<=8'd154;
		data_a[11449]<=8'd154;
		data_a[11450]<=8'd150;
		data_a[11451]<=8'd161;
		data_a[11452]<=8'd159;
		data_a[11453]<=8'd159;
		data_a[11454]<=8'd158;
		data_a[11455]<=8'd161;
		data_a[11456]<=8'd158;
		data_a[11457]<=8'd154;
		data_a[11458]<=8'd149;
		data_a[11459]<=8'd144;
		data_a[11460]<=8'd144;
		data_a[11461]<=8'd148;
		data_a[11462]<=8'd142;
		data_a[11463]<=8'd129;
		data_a[11464]<=8'd87;
		data_a[11465]<=8'd69;
		data_a[11466]<=8'd58;
		data_a[11467]<=8'd60;
		data_a[11468]<=8'd66;
		data_a[11469]<=8'd67;
		data_a[11470]<=8'd81;
		data_a[11471]<=8'd85;
		data_a[11472]<=8'd100;
		data_a[11473]<=8'd110;
		data_a[11474]<=8'd179;
		data_a[11475]<=8'd195;
		data_a[11476]<=8'd187;
		data_a[11477]<=8'd187;
		data_a[11478]<=8'd199;
		data_a[11479]<=8'd188;
		data_a[11480]<=8'd200;
		data_a[11481]<=8'd68;
		data_a[11482]<=8'd129;
		data_a[11483]<=8'd136;
		data_a[11484]<=8'd132;
		data_a[11485]<=8'd117;
		data_a[11486]<=8'd94;
		data_a[11487]<=8'd83;
		data_a[11488]<=8'd91;
		data_a[11489]<=8'd90;
		data_a[11490]<=8'd97;
		data_a[11491]<=8'd91;
		data_a[11492]<=8'd101;
		data_a[11493]<=8'd107;
		data_a[11494]<=8'd94;
		data_a[11495]<=8'd106;
		data_a[11496]<=8'd111;
		data_a[11497]<=8'd105;
		data_a[11498]<=8'd134;
		data_a[11499]<=8'd154;
		data_a[11500]<=8'd162;
		data_a[11501]<=8'd192;
		data_a[11502]<=8'd220;
		data_a[11503]<=8'd230;
		data_a[11504]<=8'd197;
		data_a[11505]<=8'd230;
		data_a[11506]<=8'd192;
		data_a[11507]<=8'd170;
		data_a[11508]<=8'd160;
		data_a[11509]<=8'd156;
		data_a[11510]<=8'd162;
		data_a[11511]<=8'd161;
		data_a[11512]<=8'd166;
		data_a[11513]<=8'd167;
		data_a[11514]<=8'd177;
		data_a[11515]<=8'd185;
		data_a[11516]<=8'd187;
		data_a[11517]<=8'd191;
		data_a[11518]<=8'd199;
		data_a[11519]<=8'd202;
		data_a[11520]<=8'd195;
		data_a[11521]<=8'd200;
		data_a[11522]<=8'd190;
		data_a[11523]<=8'd189;
		data_a[11524]<=8'd180;
		data_a[11525]<=8'd183;
		data_a[11526]<=8'd173;
		data_a[11527]<=8'd168;
		data_a[11528]<=8'd111;
		data_a[11529]<=8'd113;
		data_a[11530]<=8'd122;
		data_a[11531]<=8'd163;
		data_a[11532]<=8'd202;
		data_a[11533]<=8'd226;
		data_a[11534]<=8'd218;
		data_a[11535]<=8'd219;
		data_a[11536]<=8'd221;
		data_a[11537]<=8'd221;
		data_a[11538]<=8'd221;
		data_a[11539]<=8'd223;
		data_a[11540]<=8'd224;
		data_a[11541]<=8'd225;
		data_a[11542]<=8'd227;
		data_a[11543]<=8'd230;
		data_a[11544]<=8'd228;
		data_a[11545]<=8'd229;
		data_a[11546]<=8'd230;
		data_a[11547]<=8'd231;
		data_a[11548]<=8'd232;
		data_a[11549]<=8'd232;
		data_a[11550]<=8'd255;
		data_a[11551]<=8'd176;
		data_a[11552]<=8'd179;
		data_a[11553]<=8'd181;
		data_a[11554]<=8'd180;
		data_a[11555]<=8'd181;
		data_a[11556]<=8'd179;
		data_a[11557]<=8'd179;
		data_a[11558]<=8'd180;
		data_a[11559]<=8'd181;
		data_a[11560]<=8'd176;
		data_a[11561]<=8'd178;
		data_a[11562]<=8'd176;
		data_a[11563]<=8'd175;
		data_a[11564]<=8'd174;
		data_a[11565]<=8'd172;
		data_a[11566]<=8'd179;
		data_a[11567]<=8'd187;
		data_a[11568]<=8'd112;
		data_a[11569]<=8'd84;
		data_a[11570]<=8'd88;
		data_a[11571]<=8'd64;
		data_a[11572]<=8'd67;
		data_a[11573]<=8'd63;
		data_a[11574]<=8'd52;
		data_a[11575]<=8'd52;
		data_a[11576]<=8'd57;
		data_a[11577]<=8'd51;
		data_a[11578]<=8'd65;
		data_a[11579]<=8'd80;
		data_a[11580]<=8'd128;
		data_a[11581]<=8'd156;
		data_a[11582]<=8'd164;
		data_a[11583]<=8'd167;
		data_a[11584]<=8'd174;
		data_a[11585]<=8'd134;
		data_a[11586]<=8'd123;
		data_a[11587]<=8'd125;
		data_a[11588]<=8'd124;
		data_a[11589]<=8'd133;
		data_a[11590]<=8'd127;
		data_a[11591]<=8'd125;
		data_a[11592]<=8'd134;
		data_a[11593]<=8'd129;
		data_a[11594]<=8'd138;
		data_a[11595]<=8'd142;
		data_a[11596]<=8'd142;
		data_a[11597]<=8'd146;
		data_a[11598]<=8'd144;
		data_a[11599]<=8'd146;
		data_a[11600]<=8'd144;
		data_a[11601]<=8'd145;
		data_a[11602]<=8'd146;
		data_a[11603]<=8'd143;
		data_a[11604]<=8'd154;
		data_a[11605]<=8'd157;
		data_a[11606]<=8'd154;
		data_a[11607]<=8'd155;
		data_a[11608]<=8'd153;
		data_a[11609]<=8'd147;
		data_a[11610]<=8'd144;
		data_a[11611]<=8'd147;
		data_a[11612]<=8'd141;
		data_a[11613]<=8'd129;
		data_a[11614]<=8'd90;
		data_a[11615]<=8'd72;
		data_a[11616]<=8'd60;
		data_a[11617]<=8'd59;
		data_a[11618]<=8'd62;
		data_a[11619]<=8'd61;
		data_a[11620]<=8'd77;
		data_a[11621]<=8'd88;
		data_a[11622]<=8'd95;
		data_a[11623]<=8'd94;
		data_a[11624]<=8'd158;
		data_a[11625]<=8'd184;
		data_a[11626]<=8'd185;
		data_a[11627]<=8'd186;
		data_a[11628]<=8'd195;
		data_a[11629]<=8'd190;
		data_a[11630]<=8'd192;
		data_a[11631]<=8'd72;
		data_a[11632]<=8'd127;
		data_a[11633]<=8'd141;
		data_a[11634]<=8'd132;
		data_a[11635]<=8'd113;
		data_a[11636]<=8'd108;
		data_a[11637]<=8'd105;
		data_a[11638]<=8'd105;
		data_a[11639]<=8'd105;
		data_a[11640]<=8'd113;
		data_a[11641]<=8'd116;
		data_a[11642]<=8'd111;
		data_a[11643]<=8'd107;
		data_a[11644]<=8'd104;
		data_a[11645]<=8'd106;
		data_a[11646]<=8'd111;
		data_a[11647]<=8'd115;
		data_a[11648]<=8'd136;
		data_a[11649]<=8'd158;
		data_a[11650]<=8'd167;
		data_a[11651]<=8'd190;
		data_a[11652]<=8'd206;
		data_a[11653]<=8'd234;
		data_a[11654]<=8'd212;
		data_a[11655]<=8'd213;
		data_a[11656]<=8'd215;
		data_a[11657]<=8'd188;
		data_a[11658]<=8'd154;
		data_a[11659]<=8'd160;
		data_a[11660]<=8'd160;
		data_a[11661]<=8'd168;
		data_a[11662]<=8'd168;
		data_a[11663]<=8'd167;
		data_a[11664]<=8'd173;
		data_a[11665]<=8'd181;
		data_a[11666]<=8'd186;
		data_a[11667]<=8'd190;
		data_a[11668]<=8'd195;
		data_a[11669]<=8'd199;
		data_a[11670]<=8'd194;
		data_a[11671]<=8'd192;
		data_a[11672]<=8'd194;
		data_a[11673]<=8'd188;
		data_a[11674]<=8'd185;
		data_a[11675]<=8'd178;
		data_a[11676]<=8'd175;
		data_a[11677]<=8'd167;
		data_a[11678]<=8'd113;
		data_a[11679]<=8'd102;
		data_a[11680]<=8'd112;
		data_a[11681]<=8'd150;
		data_a[11682]<=8'd196;
		data_a[11683]<=8'd215;
		data_a[11684]<=8'd226;
		data_a[11685]<=8'd220;
		data_a[11686]<=8'd221;
		data_a[11687]<=8'd221;
		data_a[11688]<=8'd223;
		data_a[11689]<=8'd226;
		data_a[11690]<=8'd227;
		data_a[11691]<=8'd227;
		data_a[11692]<=8'd228;
		data_a[11693]<=8'd230;
		data_a[11694]<=8'd229;
		data_a[11695]<=8'd229;
		data_a[11696]<=8'd230;
		data_a[11697]<=8'd231;
		data_a[11698]<=8'd232;
		data_a[11699]<=8'd232;
		data_a[11700]<=8'd255;
		data_a[11701]<=8'd171;
		data_a[11702]<=8'd175;
		data_a[11703]<=8'd179;
		data_a[11704]<=8'd178;
		data_a[11705]<=8'd178;
		data_a[11706]<=8'd175;
		data_a[11707]<=8'd177;
		data_a[11708]<=8'd176;
		data_a[11709]<=8'd181;
		data_a[11710]<=8'd180;
		data_a[11711]<=8'd173;
		data_a[11712]<=8'd173;
		data_a[11713]<=8'd173;
		data_a[11714]<=8'd168;
		data_a[11715]<=8'd177;
		data_a[11716]<=8'd175;
		data_a[11717]<=8'd165;
		data_a[11718]<=8'd127;
		data_a[11719]<=8'd62;
		data_a[11720]<=8'd66;
		data_a[11721]<=8'd67;
		data_a[11722]<=8'd61;
		data_a[11723]<=8'd57;
		data_a[11724]<=8'd58;
		data_a[11725]<=8'd52;
		data_a[11726]<=8'd55;
		data_a[11727]<=8'd53;
		data_a[11728]<=8'd64;
		data_a[11729]<=8'd84;
		data_a[11730]<=8'd131;
		data_a[11731]<=8'd152;
		data_a[11732]<=8'd172;
		data_a[11733]<=8'd151;
		data_a[11734]<=8'd82;
		data_a[11735]<=8'd80;
		data_a[11736]<=8'd75;
		data_a[11737]<=8'd77;
		data_a[11738]<=8'd67;
		data_a[11739]<=8'd72;
		data_a[11740]<=8'd81;
		data_a[11741]<=8'd84;
		data_a[11742]<=8'd101;
		data_a[11743]<=8'd115;
		data_a[11744]<=8'd122;
		data_a[11745]<=8'd133;
		data_a[11746]<=8'd141;
		data_a[11747]<=8'd138;
		data_a[11748]<=8'd135;
		data_a[11749]<=8'd137;
		data_a[11750]<=8'd132;
		data_a[11751]<=8'd135;
		data_a[11752]<=8'd132;
		data_a[11753]<=8'd139;
		data_a[11754]<=8'd138;
		data_a[11755]<=8'd138;
		data_a[11756]<=8'd143;
		data_a[11757]<=8'd152;
		data_a[11758]<=8'd157;
		data_a[11759]<=8'd151;
		data_a[11760]<=8'd146;
		data_a[11761]<=8'd146;
		data_a[11762]<=8'd142;
		data_a[11763]<=8'd132;
		data_a[11764]<=8'd85;
		data_a[11765]<=8'd64;
		data_a[11766]<=8'd60;
		data_a[11767]<=8'd56;
		data_a[11768]<=8'd60;
		data_a[11769]<=8'd65;
		data_a[11770]<=8'd78;
		data_a[11771]<=8'd100;
		data_a[11772]<=8'd100;
		data_a[11773]<=8'd92;
		data_a[11774]<=8'd186;
		data_a[11775]<=8'd185;
		data_a[11776]<=8'd189;
		data_a[11777]<=8'd186;
		data_a[11778]<=8'd181;
		data_a[11779]<=8'd187;
		data_a[11780]<=8'd199;
		data_a[11781]<=8'd77;
		data_a[11782]<=8'd121;
		data_a[11783]<=8'd139;
		data_a[11784]<=8'd132;
		data_a[11785]<=8'd118;
		data_a[11786]<=8'd113;
		data_a[11787]<=8'd126;
		data_a[11788]<=8'd113;
		data_a[11789]<=8'd116;
		data_a[11790]<=8'd117;
		data_a[11791]<=8'd107;
		data_a[11792]<=8'd107;
		data_a[11793]<=8'd108;
		data_a[11794]<=8'd114;
		data_a[11795]<=8'd112;
		data_a[11796]<=8'd113;
		data_a[11797]<=8'd127;
		data_a[11798]<=8'd143;
		data_a[11799]<=8'd160;
		data_a[11800]<=8'd160;
		data_a[11801]<=8'd189;
		data_a[11802]<=8'd205;
		data_a[11803]<=8'd207;
		data_a[11804]<=8'd205;
		data_a[11805]<=8'd223;
		data_a[11806]<=8'd207;
		data_a[11807]<=8'd198;
		data_a[11808]<=8'd179;
		data_a[11809]<=8'd155;
		data_a[11810]<=8'd160;
		data_a[11811]<=8'd163;
		data_a[11812]<=8'd168;
		data_a[11813]<=8'd168;
		data_a[11814]<=8'd171;
		data_a[11815]<=8'd180;
		data_a[11816]<=8'd191;
		data_a[11817]<=8'd194;
		data_a[11818]<=8'd195;
		data_a[11819]<=8'd198;
		data_a[11820]<=8'd196;
		data_a[11821]<=8'd184;
		data_a[11822]<=8'd185;
		data_a[11823]<=8'd196;
		data_a[11824]<=8'd179;
		data_a[11825]<=8'd178;
		data_a[11826]<=8'd171;
		data_a[11827]<=8'd167;
		data_a[11828]<=8'd108;
		data_a[11829]<=8'd110;
		data_a[11830]<=8'd101;
		data_a[11831]<=8'd149;
		data_a[11832]<=8'd180;
		data_a[11833]<=8'd222;
		data_a[11834]<=8'd219;
		data_a[11835]<=8'd225;
		data_a[11836]<=8'd222;
		data_a[11837]<=8'd222;
		data_a[11838]<=8'd224;
		data_a[11839]<=8'd227;
		data_a[11840]<=8'd228;
		data_a[11841]<=8'd228;
		data_a[11842]<=8'd229;
		data_a[11843]<=8'd231;
		data_a[11844]<=8'd233;
		data_a[11845]<=8'd233;
		data_a[11846]<=8'd234;
		data_a[11847]<=8'd234;
		data_a[11848]<=8'd235;
		data_a[11849]<=8'd234;
		data_a[11850]<=8'd254;
		data_a[11851]<=8'd171;
		data_a[11852]<=8'd175;
		data_a[11853]<=8'd173;
		data_a[11854]<=8'd174;
		data_a[11855]<=8'd182;
		data_a[11856]<=8'd179;
		data_a[11857]<=8'd174;
		data_a[11858]<=8'd179;
		data_a[11859]<=8'd174;
		data_a[11860]<=8'd173;
		data_a[11861]<=8'd171;
		data_a[11862]<=8'd178;
		data_a[11863]<=8'd167;
		data_a[11864]<=8'd164;
		data_a[11865]<=8'd159;
		data_a[11866]<=8'd163;
		data_a[11867]<=8'd181;
		data_a[11868]<=8'd182;
		data_a[11869]<=8'd71;
		data_a[11870]<=8'd68;
		data_a[11871]<=8'd65;
		data_a[11872]<=8'd53;
		data_a[11873]<=8'd60;
		data_a[11874]<=8'd61;
		data_a[11875]<=8'd50;
		data_a[11876]<=8'd55;
		data_a[11877]<=8'd54;
		data_a[11878]<=8'd60;
		data_a[11879]<=8'd84;
		data_a[11880]<=8'd132;
		data_a[11881]<=8'd147;
		data_a[11882]<=8'd115;
		data_a[11883]<=8'd89;
		data_a[11884]<=8'd80;
		data_a[11885]<=8'd79;
		data_a[11886]<=8'd67;
		data_a[11887]<=8'd67;
		data_a[11888]<=8'd63;
		data_a[11889]<=8'd62;
		data_a[11890]<=8'd62;
		data_a[11891]<=8'd73;
		data_a[11892]<=8'd73;
		data_a[11893]<=8'd91;
		data_a[11894]<=8'd106;
		data_a[11895]<=8'd122;
		data_a[11896]<=8'd130;
		data_a[11897]<=8'd135;
		data_a[11898]<=8'd128;
		data_a[11899]<=8'd125;
		data_a[11900]<=8'd121;
		data_a[11901]<=8'd114;
		data_a[11902]<=8'd111;
		data_a[11903]<=8'd120;
		data_a[11904]<=8'd121;
		data_a[11905]<=8'd127;
		data_a[11906]<=8'd132;
		data_a[11907]<=8'd147;
		data_a[11908]<=8'd158;
		data_a[11909]<=8'd153;
		data_a[11910]<=8'd145;
		data_a[11911]<=8'd144;
		data_a[11912]<=8'd142;
		data_a[11913]<=8'd134;
		data_a[11914]<=8'd91;
		data_a[11915]<=8'd62;
		data_a[11916]<=8'd62;
		data_a[11917]<=8'd55;
		data_a[11918]<=8'd62;
		data_a[11919]<=8'd68;
		data_a[11920]<=8'd68;
		data_a[11921]<=8'd88;
		data_a[11922]<=8'd92;
		data_a[11923]<=8'd110;
		data_a[11924]<=8'd176;
		data_a[11925]<=8'd184;
		data_a[11926]<=8'd179;
		data_a[11927]<=8'd187;
		data_a[11928]<=8'd178;
		data_a[11929]<=8'd184;
		data_a[11930]<=8'd164;
		data_a[11931]<=8'd78;
		data_a[11932]<=8'd120;
		data_a[11933]<=8'd144;
		data_a[11934]<=8'd142;
		data_a[11935]<=8'd134;
		data_a[11936]<=8'd136;
		data_a[11937]<=8'd135;
		data_a[11938]<=8'd117;
		data_a[11939]<=8'd119;
		data_a[11940]<=8'd111;
		data_a[11941]<=8'd109;
		data_a[11942]<=8'd119;
		data_a[11943]<=8'd117;
		data_a[11944]<=8'd119;
		data_a[11945]<=8'd119;
		data_a[11946]<=8'd128;
		data_a[11947]<=8'd141;
		data_a[11948]<=8'd144;
		data_a[11949]<=8'd157;
		data_a[11950]<=8'd169;
		data_a[11951]<=8'd184;
		data_a[11952]<=8'd201;
		data_a[11953]<=8'd198;
		data_a[11954]<=8'd196;
		data_a[11955]<=8'd206;
		data_a[11956]<=8'd221;
		data_a[11957]<=8'd194;
		data_a[11958]<=8'd198;
		data_a[11959]<=8'd198;
		data_a[11960]<=8'd154;
		data_a[11961]<=8'd158;
		data_a[11962]<=8'd157;
		data_a[11963]<=8'd162;
		data_a[11964]<=8'd168;
		data_a[11965]<=8'd176;
		data_a[11966]<=8'd185;
		data_a[11967]<=8'd185;
		data_a[11968]<=8'd185;
		data_a[11969]<=8'd191;
		data_a[11970]<=8'd189;
		data_a[11971]<=8'd185;
		data_a[11972]<=8'd182;
		data_a[11973]<=8'd184;
		data_a[11974]<=8'd180;
		data_a[11975]<=8'd177;
		data_a[11976]<=8'd168;
		data_a[11977]<=8'd166;
		data_a[11978]<=8'd103;
		data_a[11979]<=8'd102;
		data_a[11980]<=8'd103;
		data_a[11981]<=8'd136;
		data_a[11982]<=8'd168;
		data_a[11983]<=8'd226;
		data_a[11984]<=8'd224;
		data_a[11985]<=8'd224;
		data_a[11986]<=8'd225;
		data_a[11987]<=8'd224;
		data_a[11988]<=8'd225;
		data_a[11989]<=8'd227;
		data_a[11990]<=8'd228;
		data_a[11991]<=8'd228;
		data_a[11992]<=8'd230;
		data_a[11993]<=8'd234;
		data_a[11994]<=8'd232;
		data_a[11995]<=8'd232;
		data_a[11996]<=8'd233;
		data_a[11997]<=8'd234;
		data_a[11998]<=8'd235;
		data_a[11999]<=8'd235;
		data_a[12000]<=8'd253;
		data_a[12001]<=8'd168;
		data_a[12002]<=8'd172;
		data_a[12003]<=8'd174;
		data_a[12004]<=8'd175;
		data_a[12005]<=8'd175;
		data_a[12006]<=8'd171;
		data_a[12007]<=8'd170;
		data_a[12008]<=8'd169;
		data_a[12009]<=8'd178;
		data_a[12010]<=8'd171;
		data_a[12011]<=8'd161;
		data_a[12012]<=8'd158;
		data_a[12013]<=8'd166;
		data_a[12014]<=8'd168;
		data_a[12015]<=8'd171;
		data_a[12016]<=8'd169;
		data_a[12017]<=8'd174;
		data_a[12018]<=8'd177;
		data_a[12019]<=8'd140;
		data_a[12020]<=8'd75;
		data_a[12021]<=8'd66;
		data_a[12022]<=8'd56;
		data_a[12023]<=8'd53;
		data_a[12024]<=8'd56;
		data_a[12025]<=8'd54;
		data_a[12026]<=8'd51;
		data_a[12027]<=8'd48;
		data_a[12028]<=8'd64;
		data_a[12029]<=8'd87;
		data_a[12030]<=8'd139;
		data_a[12031]<=8'd143;
		data_a[12032]<=8'd98;
		data_a[12033]<=8'd101;
		data_a[12034]<=8'd104;
		data_a[12035]<=8'd109;
		data_a[12036]<=8'd95;
		data_a[12037]<=8'd81;
		data_a[12038]<=8'd73;
		data_a[12039]<=8'd63;
		data_a[12040]<=8'd58;
		data_a[12041]<=8'd60;
		data_a[12042]<=8'd70;
		data_a[12043]<=8'd73;
		data_a[12044]<=8'd98;
		data_a[12045]<=8'd113;
		data_a[12046]<=8'd124;
		data_a[12047]<=8'd124;
		data_a[12048]<=8'd125;
		data_a[12049]<=8'd119;
		data_a[12050]<=8'd108;
		data_a[12051]<=8'd97;
		data_a[12052]<=8'd90;
		data_a[12053]<=8'd88;
		data_a[12054]<=8'd90;
		data_a[12055]<=8'd98;
		data_a[12056]<=8'd105;
		data_a[12057]<=8'd119;
		data_a[12058]<=8'd134;
		data_a[12059]<=8'd153;
		data_a[12060]<=8'd152;
		data_a[12061]<=8'd146;
		data_a[12062]<=8'd140;
		data_a[12063]<=8'd134;
		data_a[12064]<=8'd85;
		data_a[12065]<=8'd60;
		data_a[12066]<=8'd56;
		data_a[12067]<=8'd58;
		data_a[12068]<=8'd58;
		data_a[12069]<=8'd60;
		data_a[12070]<=8'd67;
		data_a[12071]<=8'd82;
		data_a[12072]<=8'd90;
		data_a[12073]<=8'd125;
		data_a[12074]<=8'd159;
		data_a[12075]<=8'd179;
		data_a[12076]<=8'd183;
		data_a[12077]<=8'd166;
		data_a[12078]<=8'd168;
		data_a[12079]<=8'd164;
		data_a[12080]<=8'd168;
		data_a[12081]<=8'd99;
		data_a[12082]<=8'd121;
		data_a[12083]<=8'd146;
		data_a[12084]<=8'd146;
		data_a[12085]<=8'd146;
		data_a[12086]<=8'd149;
		data_a[12087]<=8'd144;
		data_a[12088]<=8'd132;
		data_a[12089]<=8'd122;
		data_a[12090]<=8'd125;
		data_a[12091]<=8'd125;
		data_a[12092]<=8'd131;
		data_a[12093]<=8'd128;
		data_a[12094]<=8'd126;
		data_a[12095]<=8'd130;
		data_a[12096]<=8'd144;
		data_a[12097]<=8'd142;
		data_a[12098]<=8'd153;
		data_a[12099]<=8'd159;
		data_a[12100]<=8'd173;
		data_a[12101]<=8'd192;
		data_a[12102]<=8'd190;
		data_a[12103]<=8'd184;
		data_a[12104]<=8'd184;
		data_a[12105]<=8'd190;
		data_a[12106]<=8'd183;
		data_a[12107]<=8'd181;
		data_a[12108]<=8'd185;
		data_a[12109]<=8'd202;
		data_a[12110]<=8'd187;
		data_a[12111]<=8'd140;
		data_a[12112]<=8'd149;
		data_a[12113]<=8'd154;
		data_a[12114]<=8'd166;
		data_a[12115]<=8'd169;
		data_a[12116]<=8'd180;
		data_a[12117]<=8'd180;
		data_a[12118]<=8'd186;
		data_a[12119]<=8'd185;
		data_a[12120]<=8'd187;
		data_a[12121]<=8'd181;
		data_a[12122]<=8'd188;
		data_a[12123]<=8'd181;
		data_a[12124]<=8'd179;
		data_a[12125]<=8'd172;
		data_a[12126]<=8'd172;
		data_a[12127]<=8'd168;
		data_a[12128]<=8'd110;
		data_a[12129]<=8'd101;
		data_a[12130]<=8'd107;
		data_a[12131]<=8'd129;
		data_a[12132]<=8'd151;
		data_a[12133]<=8'd200;
		data_a[12134]<=8'd228;
		data_a[12135]<=8'd226;
		data_a[12136]<=8'd228;
		data_a[12137]<=8'd227;
		data_a[12138]<=8'd227;
		data_a[12139]<=8'd228;
		data_a[12140]<=8'd230;
		data_a[12141]<=8'd232;
		data_a[12142]<=8'd232;
		data_a[12143]<=8'd232;
		data_a[12144]<=8'd234;
		data_a[12145]<=8'd235;
		data_a[12146]<=8'd235;
		data_a[12147]<=8'd235;
		data_a[12148]<=8'd235;
		data_a[12149]<=8'd236;
		data_a[12150]<=8'd255;
		data_a[12151]<=8'd146;
		data_a[12152]<=8'd160;
		data_a[12153]<=8'd168;
		data_a[12154]<=8'd175;
		data_a[12155]<=8'd162;
		data_a[12156]<=8'd180;
		data_a[12157]<=8'd167;
		data_a[12158]<=8'd151;
		data_a[12159]<=8'd158;
		data_a[12160]<=8'd166;
		data_a[12161]<=8'd163;
		data_a[12162]<=8'd174;
		data_a[12163]<=8'd170;
		data_a[12164]<=8'd162;
		data_a[12165]<=8'd171;
		data_a[12166]<=8'd166;
		data_a[12167]<=8'd164;
		data_a[12168]<=8'd167;
		data_a[12169]<=8'd175;
		data_a[12170]<=8'd74;
		data_a[12171]<=8'd64;
		data_a[12172]<=8'd55;
		data_a[12173]<=8'd56;
		data_a[12174]<=8'd55;
		data_a[12175]<=8'd59;
		data_a[12176]<=8'd51;
		data_a[12177]<=8'd53;
		data_a[12178]<=8'd49;
		data_a[12179]<=8'd106;
		data_a[12180]<=8'd57;
		data_a[12181]<=8'd51;
		data_a[12182]<=8'd68;
		data_a[12183]<=8'd57;
		data_a[12184]<=8'd61;
		data_a[12185]<=8'd69;
		data_a[12186]<=8'd64;
		data_a[12187]<=8'd66;
		data_a[12188]<=8'd74;
		data_a[12189]<=8'd78;
		data_a[12190]<=8'd64;
		data_a[12191]<=8'd66;
		data_a[12192]<=8'd70;
		data_a[12193]<=8'd66;
		data_a[12194]<=8'd82;
		data_a[12195]<=8'd105;
		data_a[12196]<=8'd110;
		data_a[12197]<=8'd119;
		data_a[12198]<=8'd105;
		data_a[12199]<=8'd115;
		data_a[12200]<=8'd94;
		data_a[12201]<=8'd87;
		data_a[12202]<=8'd69;
		data_a[12203]<=8'd66;
		data_a[12204]<=8'd68;
		data_a[12205]<=8'd63;
		data_a[12206]<=8'd67;
		data_a[12207]<=8'd76;
		data_a[12208]<=8'd80;
		data_a[12209]<=8'd110;
		data_a[12210]<=8'd141;
		data_a[12211]<=8'd146;
		data_a[12212]<=8'd144;
		data_a[12213]<=8'd130;
		data_a[12214]<=8'd82;
		data_a[12215]<=8'd66;
		data_a[12216]<=8'd59;
		data_a[12217]<=8'd52;
		data_a[12218]<=8'd57;
		data_a[12219]<=8'd63;
		data_a[12220]<=8'd68;
		data_a[12221]<=8'd78;
		data_a[12222]<=8'd98;
		data_a[12223]<=8'd131;
		data_a[12224]<=8'd144;
		data_a[12225]<=8'd172;
		data_a[12226]<=8'd159;
		data_a[12227]<=8'd181;
		data_a[12228]<=8'd182;
		data_a[12229]<=8'd182;
		data_a[12230]<=8'd180;
		data_a[12231]<=8'd117;
		data_a[12232]<=8'd128;
		data_a[12233]<=8'd146;
		data_a[12234]<=8'd149;
		data_a[12235]<=8'd157;
		data_a[12236]<=8'd152;
		data_a[12237]<=8'd150;
		data_a[12238]<=8'd152;
		data_a[12239]<=8'd145;
		data_a[12240]<=8'd138;
		data_a[12241]<=8'd134;
		data_a[12242]<=8'd129;
		data_a[12243]<=8'd135;
		data_a[12244]<=8'd137;
		data_a[12245]<=8'd146;
		data_a[12246]<=8'd148;
		data_a[12247]<=8'd152;
		data_a[12248]<=8'd144;
		data_a[12249]<=8'd153;
		data_a[12250]<=8'd180;
		data_a[12251]<=8'd189;
		data_a[12252]<=8'd181;
		data_a[12253]<=8'd172;
		data_a[12254]<=8'd166;
		data_a[12255]<=8'd163;
		data_a[12256]<=8'd164;
		data_a[12257]<=8'd160;
		data_a[12258]<=8'd164;
		data_a[12259]<=8'd165;
		data_a[12260]<=8'd179;
		data_a[12261]<=8'd158;
		data_a[12262]<=8'd141;
		data_a[12263]<=8'd145;
		data_a[12264]<=8'd154;
		data_a[12265]<=8'd165;
		data_a[12266]<=8'd170;
		data_a[12267]<=8'd176;
		data_a[12268]<=8'd177;
		data_a[12269]<=8'd182;
		data_a[12270]<=8'd184;
		data_a[12271]<=8'd182;
		data_a[12272]<=8'd179;
		data_a[12273]<=8'd182;
		data_a[12274]<=8'd173;
		data_a[12275]<=8'd165;
		data_a[12276]<=8'd167;
		data_a[12277]<=8'd166;
		data_a[12278]<=8'd106;
		data_a[12279]<=8'd103;
		data_a[12280]<=8'd109;
		data_a[12281]<=8'd127;
		data_a[12282]<=8'd160;
		data_a[12283]<=8'd193;
		data_a[12284]<=8'd222;
		data_a[12285]<=8'd225;
		data_a[12286]<=8'd228;
		data_a[12287]<=8'd227;
		data_a[12288]<=8'd227;
		data_a[12289]<=8'd229;
		data_a[12290]<=8'd231;
		data_a[12291]<=8'd233;
		data_a[12292]<=8'd233;
		data_a[12293]<=8'd233;
		data_a[12294]<=8'd234;
		data_a[12295]<=8'd236;
		data_a[12296]<=8'd236;
		data_a[12297]<=8'd236;
		data_a[12298]<=8'd237;
		data_a[12299]<=8'd238;
		data_a[12300]<=8'd254;
		data_a[12301]<=8'd150;
		data_a[12302]<=8'd144;
		data_a[12303]<=8'd150;
		data_a[12304]<=8'd145;
		data_a[12305]<=8'd159;
		data_a[12306]<=8'd159;
		data_a[12307]<=8'd172;
		data_a[12308]<=8'd172;
		data_a[12309]<=8'd166;
		data_a[12310]<=8'd169;
		data_a[12311]<=8'd161;
		data_a[12312]<=8'd161;
		data_a[12313]<=8'd163;
		data_a[12314]<=8'd166;
		data_a[12315]<=8'd164;
		data_a[12316]<=8'd166;
		data_a[12317]<=8'd171;
		data_a[12318]<=8'd165;
		data_a[12319]<=8'd158;
		data_a[12320]<=8'd95;
		data_a[12321]<=8'd60;
		data_a[12322]<=8'd59;
		data_a[12323]<=8'd63;
		data_a[12324]<=8'd67;
		data_a[12325]<=8'd51;
		data_a[12326]<=8'd52;
		data_a[12327]<=8'd58;
		data_a[12328]<=8'd61;
		data_a[12329]<=8'd67;
		data_a[12330]<=8'd62;
		data_a[12331]<=8'd58;
		data_a[12332]<=8'd99;
		data_a[12333]<=8'd115;
		data_a[12334]<=8'd109;
		data_a[12335]<=8'd105;
		data_a[12336]<=8'd100;
		data_a[12337]<=8'd92;
		data_a[12338]<=8'd99;
		data_a[12339]<=8'd95;
		data_a[12340]<=8'd93;
		data_a[12341]<=8'd67;
		data_a[12342]<=8'd73;
		data_a[12343]<=8'd80;
		data_a[12344]<=8'd74;
		data_a[12345]<=8'd92;
		data_a[12346]<=8'd114;
		data_a[12347]<=8'd113;
		data_a[12348]<=8'd112;
		data_a[12349]<=8'd103;
		data_a[12350]<=8'd89;
		data_a[12351]<=8'd74;
		data_a[12352]<=8'd69;
		data_a[12353]<=8'd59;
		data_a[12354]<=8'd58;
		data_a[12355]<=8'd52;
		data_a[12356]<=8'd58;
		data_a[12357]<=8'd55;
		data_a[12358]<=8'd59;
		data_a[12359]<=8'd74;
		data_a[12360]<=8'd109;
		data_a[12361]<=8'd145;
		data_a[12362]<=8'd129;
		data_a[12363]<=8'd143;
		data_a[12364]<=8'd87;
		data_a[12365]<=8'd58;
		data_a[12366]<=8'd59;
		data_a[12367]<=8'd54;
		data_a[12368]<=8'd58;
		data_a[12369]<=8'd53;
		data_a[12370]<=8'd75;
		data_a[12371]<=8'd84;
		data_a[12372]<=8'd77;
		data_a[12373]<=8'd91;
		data_a[12374]<=8'd178;
		data_a[12375]<=8'd153;
		data_a[12376]<=8'd167;
		data_a[12377]<=8'd176;
		data_a[12378]<=8'd186;
		data_a[12379]<=8'd186;
		data_a[12380]<=8'd188;
		data_a[12381]<=8'd182;
		data_a[12382]<=8'd103;
		data_a[12383]<=8'd154;
		data_a[12384]<=8'd153;
		data_a[12385]<=8'd158;
		data_a[12386]<=8'd163;
		data_a[12387]<=8'd160;
		data_a[12388]<=8'd162;
		data_a[12389]<=8'd160;
		data_a[12390]<=8'd154;
		data_a[12391]<=8'd150;
		data_a[12392]<=8'd145;
		data_a[12393]<=8'd151;
		data_a[12394]<=8'd151;
		data_a[12395]<=8'd156;
		data_a[12396]<=8'd152;
		data_a[12397]<=8'd149;
		data_a[12398]<=8'd151;
		data_a[12399]<=8'd179;
		data_a[12400]<=8'd173;
		data_a[12401]<=8'd151;
		data_a[12402]<=8'd165;
		data_a[12403]<=8'd162;
		data_a[12404]<=8'd156;
		data_a[12405]<=8'd150;
		data_a[12406]<=8'd138;
		data_a[12407]<=8'd140;
		data_a[12408]<=8'd138;
		data_a[12409]<=8'd140;
		data_a[12410]<=8'd153;
		data_a[12411]<=8'd155;
		data_a[12412]<=8'd147;
		data_a[12413]<=8'd141;
		data_a[12414]<=8'd146;
		data_a[12415]<=8'd156;
		data_a[12416]<=8'd154;
		data_a[12417]<=8'd169;
		data_a[12418]<=8'd171;
		data_a[12419]<=8'd173;
		data_a[12420]<=8'd175;
		data_a[12421]<=8'd177;
		data_a[12422]<=8'd175;
		data_a[12423]<=8'd185;
		data_a[12424]<=8'd178;
		data_a[12425]<=8'd163;
		data_a[12426]<=8'd168;
		data_a[12427]<=8'd167;
		data_a[12428]<=8'd109;
		data_a[12429]<=8'd106;
		data_a[12430]<=8'd105;
		data_a[12431]<=8'd158;
		data_a[12432]<=8'd193;
		data_a[12433]<=8'd191;
		data_a[12434]<=8'd228;
		data_a[12435]<=8'd226;
		data_a[12436]<=8'd229;
		data_a[12437]<=8'd228;
		data_a[12438]<=8'd228;
		data_a[12439]<=8'd230;
		data_a[12440]<=8'd232;
		data_a[12441]<=8'd233;
		data_a[12442]<=8'd234;
		data_a[12443]<=8'd234;
		data_a[12444]<=8'd234;
		data_a[12445]<=8'd235;
		data_a[12446]<=8'd236;
		data_a[12447]<=8'd236;
		data_a[12448]<=8'd237;
		data_a[12449]<=8'd238;
		data_a[12450]<=8'd255;
		data_a[12451]<=8'd81;
		data_a[12452]<=8'd122;
		data_a[12453]<=8'd143;
		data_a[12454]<=8'd146;
		data_a[12455]<=8'd147;
		data_a[12456]<=8'd157;
		data_a[12457]<=8'd154;
		data_a[12458]<=8'd162;
		data_a[12459]<=8'd165;
		data_a[12460]<=8'd162;
		data_a[12461]<=8'd164;
		data_a[12462]<=8'd165;
		data_a[12463]<=8'd158;
		data_a[12464]<=8'd158;
		data_a[12465]<=8'd162;
		data_a[12466]<=8'd162;
		data_a[12467]<=8'd162;
		data_a[12468]<=8'd164;
		data_a[12469]<=8'd171;
		data_a[12470]<=8'd72;
		data_a[12471]<=8'd61;
		data_a[12472]<=8'd68;
		data_a[12473]<=8'd57;
		data_a[12474]<=8'd80;
		data_a[12475]<=8'd55;
		data_a[12476]<=8'd47;
		data_a[12477]<=8'd54;
		data_a[12478]<=8'd59;
		data_a[12479]<=8'd60;
		data_a[12480]<=8'd53;
		data_a[12481]<=8'd120;
		data_a[12482]<=8'd107;
		data_a[12483]<=8'd100;
		data_a[12484]<=8'd93;
		data_a[12485]<=8'd74;
		data_a[12486]<=8'd68;
		data_a[12487]<=8'd84;
		data_a[12488]<=8'd83;
		data_a[12489]<=8'd71;
		data_a[12490]<=8'd72;
		data_a[12491]<=8'd70;
		data_a[12492]<=8'd82;
		data_a[12493]<=8'd99;
		data_a[12494]<=8'd67;
		data_a[12495]<=8'd63;
		data_a[12496]<=8'd87;
		data_a[12497]<=8'd93;
		data_a[12498]<=8'd85;
		data_a[12499]<=8'd84;
		data_a[12500]<=8'd78;
		data_a[12501]<=8'd89;
		data_a[12502]<=8'd73;
		data_a[12503]<=8'd51;
		data_a[12504]<=8'd54;
		data_a[12505]<=8'd61;
		data_a[12506]<=8'd53;
		data_a[12507]<=8'd54;
		data_a[12508]<=8'd50;
		data_a[12509]<=8'd52;
		data_a[12510]<=8'd67;
		data_a[12511]<=8'd78;
		data_a[12512]<=8'd129;
		data_a[12513]<=8'd133;
		data_a[12514]<=8'd91;
		data_a[12515]<=8'd63;
		data_a[12516]<=8'd55;
		data_a[12517]<=8'd54;
		data_a[12518]<=8'd65;
		data_a[12519]<=8'd61;
		data_a[12520]<=8'd67;
		data_a[12521]<=8'd95;
		data_a[12522]<=8'd142;
		data_a[12523]<=8'd175;
		data_a[12524]<=8'd171;
		data_a[12525]<=8'd175;
		data_a[12526]<=8'd178;
		data_a[12527]<=8'd196;
		data_a[12528]<=8'd195;
		data_a[12529]<=8'd195;
		data_a[12530]<=8'd199;
		data_a[12531]<=8'd210;
		data_a[12532]<=8'd97;
		data_a[12533]<=8'd147;
		data_a[12534]<=8'd157;
		data_a[12535]<=8'd158;
		data_a[12536]<=8'd165;
		data_a[12537]<=8'd170;
		data_a[12538]<=8'd170;
		data_a[12539]<=8'd165;
		data_a[12540]<=8'd164;
		data_a[12541]<=8'd158;
		data_a[12542]<=8'd163;
		data_a[12543]<=8'd163;
		data_a[12544]<=8'd165;
		data_a[12545]<=8'd162;
		data_a[12546]<=8'd165;
		data_a[12547]<=8'd150;
		data_a[12548]<=8'd181;
		data_a[12549]<=8'd177;
		data_a[12550]<=8'd140;
		data_a[12551]<=8'd139;
		data_a[12552]<=8'd145;
		data_a[12553]<=8'd142;
		data_a[12554]<=8'd132;
		data_a[12555]<=8'd133;
		data_a[12556]<=8'd121;
		data_a[12557]<=8'd109;
		data_a[12558]<=8'd60;
		data_a[12559]<=8'd100;
		data_a[12560]<=8'd128;
		data_a[12561]<=8'd142;
		data_a[12562]<=8'd156;
		data_a[12563]<=8'd148;
		data_a[12564]<=8'd142;
		data_a[12565]<=8'd131;
		data_a[12566]<=8'd139;
		data_a[12567]<=8'd153;
		data_a[12568]<=8'd157;
		data_a[12569]<=8'd160;
		data_a[12570]<=8'd167;
		data_a[12571]<=8'd168;
		data_a[12572]<=8'd173;
		data_a[12573]<=8'd176;
		data_a[12574]<=8'd176;
		data_a[12575]<=8'd157;
		data_a[12576]<=8'd160;
		data_a[12577]<=8'd157;
		data_a[12578]<=8'd112;
		data_a[12579]<=8'd92;
		data_a[12580]<=8'd99;
		data_a[12581]<=8'd170;
		data_a[12582]<=8'd196;
		data_a[12583]<=8'd189;
		data_a[12584]<=8'd224;
		data_a[12585]<=8'd231;
		data_a[12586]<=8'd229;
		data_a[12587]<=8'd229;
		data_a[12588]<=8'd230;
		data_a[12589]<=8'd231;
		data_a[12590]<=8'd232;
		data_a[12591]<=8'd233;
		data_a[12592]<=8'd234;
		data_a[12593]<=8'd235;
		data_a[12594]<=8'd234;
		data_a[12595]<=8'd236;
		data_a[12596]<=8'd236;
		data_a[12597]<=8'd237;
		data_a[12598]<=8'd237;
		data_a[12599]<=8'd239;
		data_a[12600]<=8'd254;
		data_a[12601]<=8'd87;
		data_a[12602]<=8'd88;
		data_a[12603]<=8'd82;
		data_a[12604]<=8'd100;
		data_a[12605]<=8'd146;
		data_a[12606]<=8'd150;
		data_a[12607]<=8'd147;
		data_a[12608]<=8'd140;
		data_a[12609]<=8'd144;
		data_a[12610]<=8'd153;
		data_a[12611]<=8'd154;
		data_a[12612]<=8'd157;
		data_a[12613]<=8'd158;
		data_a[12614]<=8'd159;
		data_a[12615]<=8'd159;
		data_a[12616]<=8'd164;
		data_a[12617]<=8'd158;
		data_a[12618]<=8'd163;
		data_a[12619]<=8'd155;
		data_a[12620]<=8'd77;
		data_a[12621]<=8'd57;
		data_a[12622]<=8'd62;
		data_a[12623]<=8'd65;
		data_a[12624]<=8'd63;
		data_a[12625]<=8'd65;
		data_a[12626]<=8'd54;
		data_a[12627]<=8'd64;
		data_a[12628]<=8'd65;
		data_a[12629]<=8'd57;
		data_a[12630]<=8'd56;
		data_a[12631]<=8'd101;
		data_a[12632]<=8'd99;
		data_a[12633]<=8'd91;
		data_a[12634]<=8'd70;
		data_a[12635]<=8'd77;
		data_a[12636]<=8'd84;
		data_a[12637]<=8'd75;
		data_a[12638]<=8'd61;
		data_a[12639]<=8'd64;
		data_a[12640]<=8'd65;
		data_a[12641]<=8'd62;
		data_a[12642]<=8'd75;
		data_a[12643]<=8'd87;
		data_a[12644]<=8'd131;
		data_a[12645]<=8'd71;
		data_a[12646]<=8'd51;
		data_a[12647]<=8'd54;
		data_a[12648]<=8'd67;
		data_a[12649]<=8'd40;
		data_a[12650]<=8'd65;
		data_a[12651]<=8'd67;
		data_a[12652]<=8'd94;
		data_a[12653]<=8'd88;
		data_a[12654]<=8'd84;
		data_a[12655]<=8'd87;
		data_a[12656]<=8'd86;
		data_a[12657]<=8'd92;
		data_a[12658]<=8'd97;
		data_a[12659]<=8'd92;
		data_a[12660]<=8'd94;
		data_a[12661]<=8'd71;
		data_a[12662]<=8'd47;
		data_a[12663]<=8'd52;
		data_a[12664]<=8'd70;
		data_a[12665]<=8'd112;
		data_a[12666]<=8'd59;
		data_a[12667]<=8'd48;
		data_a[12668]<=8'd54;
		data_a[12669]<=8'd54;
		data_a[12670]<=8'd77;
		data_a[12671]<=8'd126;
		data_a[12672]<=8'd164;
		data_a[12673]<=8'd178;
		data_a[12674]<=8'd180;
		data_a[12675]<=8'd186;
		data_a[12676]<=8'd174;
		data_a[12677]<=8'd199;
		data_a[12678]<=8'd199;
		data_a[12679]<=8'd201;
		data_a[12680]<=8'd203;
		data_a[12681]<=8'd204;
		data_a[12682]<=8'd95;
		data_a[12683]<=8'd148;
		data_a[12684]<=8'd152;
		data_a[12685]<=8'd164;
		data_a[12686]<=8'd164;
		data_a[12687]<=8'd171;
		data_a[12688]<=8'd173;
		data_a[12689]<=8'd171;
		data_a[12690]<=8'd172;
		data_a[12691]<=8'd171;
		data_a[12692]<=8'd177;
		data_a[12693]<=8'd173;
		data_a[12694]<=8'd171;
		data_a[12695]<=8'd164;
		data_a[12696]<=8'd160;
		data_a[12697]<=8'd157;
		data_a[12698]<=8'd168;
		data_a[12699]<=8'd161;
		data_a[12700]<=8'd135;
		data_a[12701]<=8'd125;
		data_a[12702]<=8'd129;
		data_a[12703]<=8'd128;
		data_a[12704]<=8'd114;
		data_a[12705]<=8'd118;
		data_a[12706]<=8'd121;
		data_a[12707]<=8'd55;
		data_a[12708]<=8'd61;
		data_a[12709]<=8'd82;
		data_a[12710]<=8'd119;
		data_a[12711]<=8'd138;
		data_a[12712]<=8'd167;
		data_a[12713]<=8'd171;
		data_a[12714]<=8'd155;
		data_a[12715]<=8'd126;
		data_a[12716]<=8'd136;
		data_a[12717]<=8'd146;
		data_a[12718]<=8'd149;
		data_a[12719]<=8'd160;
		data_a[12720]<=8'd160;
		data_a[12721]<=8'd160;
		data_a[12722]<=8'd168;
		data_a[12723]<=8'd163;
		data_a[12724]<=8'd166;
		data_a[12725]<=8'd157;
		data_a[12726]<=8'd156;
		data_a[12727]<=8'd154;
		data_a[12728]<=8'd100;
		data_a[12729]<=8'd98;
		data_a[12730]<=8'd103;
		data_a[12731]<=8'd178;
		data_a[12732]<=8'd212;
		data_a[12733]<=8'd191;
		data_a[12734]<=8'd235;
		data_a[12735]<=8'd225;
		data_a[12736]<=8'd230;
		data_a[12737]<=8'd231;
		data_a[12738]<=8'd231;
		data_a[12739]<=8'd232;
		data_a[12740]<=8'd232;
		data_a[12741]<=8'd233;
		data_a[12742]<=8'd234;
		data_a[12743]<=8'd235;
		data_a[12744]<=8'd236;
		data_a[12745]<=8'd237;
		data_a[12746]<=8'd238;
		data_a[12747]<=8'd238;
		data_a[12748]<=8'd239;
		data_a[12749]<=8'd241;
		data_a[12750]<=8'd255;
		data_a[12751]<=8'd93;
		data_a[12752]<=8'd88;
		data_a[12753]<=8'd87;
		data_a[12754]<=8'd87;
		data_a[12755]<=8'd79;
		data_a[12756]<=8'd100;
		data_a[12757]<=8'd142;
		data_a[12758]<=8'd148;
		data_a[12759]<=8'd141;
		data_a[12760]<=8'd146;
		data_a[12761]<=8'd141;
		data_a[12762]<=8'd157;
		data_a[12763]<=8'd165;
		data_a[12764]<=8'd155;
		data_a[12765]<=8'd160;
		data_a[12766]<=8'd159;
		data_a[12767]<=8'd150;
		data_a[12768]<=8'd147;
		data_a[12769]<=8'd144;
		data_a[12770]<=8'd60;
		data_a[12771]<=8'd59;
		data_a[12772]<=8'd54;
		data_a[12773]<=8'd58;
		data_a[12774]<=8'd66;
		data_a[12775]<=8'd72;
		data_a[12776]<=8'd58;
		data_a[12777]<=8'd63;
		data_a[12778]<=8'd66;
		data_a[12779]<=8'd82;
		data_a[12780]<=8'd60;
		data_a[12781]<=8'd108;
		data_a[12782]<=8'd93;
		data_a[12783]<=8'd85;
		data_a[12784]<=8'd79;
		data_a[12785]<=8'd64;
		data_a[12786]<=8'd60;
		data_a[12787]<=8'd84;
		data_a[12788]<=8'd61;
		data_a[12789]<=8'd59;
		data_a[12790]<=8'd65;
		data_a[12791]<=8'd64;
		data_a[12792]<=8'd77;
		data_a[12793]<=8'd96;
		data_a[12794]<=8'd98;
		data_a[12795]<=8'd59;
		data_a[12796]<=8'd48;
		data_a[12797]<=8'd73;
		data_a[12798]<=8'd42;
		data_a[12799]<=8'd48;
		data_a[12800]<=8'd77;
		data_a[12801]<=8'd82;
		data_a[12802]<=8'd87;
		data_a[12803]<=8'd87;
		data_a[12804]<=8'd81;
		data_a[12805]<=8'd74;
		data_a[12806]<=8'd82;
		data_a[12807]<=8'd85;
		data_a[12808]<=8'd93;
		data_a[12809]<=8'd97;
		data_a[12810]<=8'd98;
		data_a[12811]<=8'd89;
		data_a[12812]<=8'd117;
		data_a[12813]<=8'd52;
		data_a[12814]<=8'd52;
		data_a[12815]<=8'd43;
		data_a[12816]<=8'd53;
		data_a[12817]<=8'd60;
		data_a[12818]<=8'd54;
		data_a[12819]<=8'd60;
		data_a[12820]<=8'd76;
		data_a[12821]<=8'd120;
		data_a[12822]<=8'd178;
		data_a[12823]<=8'd180;
		data_a[12824]<=8'd188;
		data_a[12825]<=8'd183;
		data_a[12826]<=8'd188;
		data_a[12827]<=8'd203;
		data_a[12828]<=8'd205;
		data_a[12829]<=8'd203;
		data_a[12830]<=8'd204;
		data_a[12831]<=8'd213;
		data_a[12832]<=8'd80;
		data_a[12833]<=8'd149;
		data_a[12834]<=8'd149;
		data_a[12835]<=8'd160;
		data_a[12836]<=8'd166;
		data_a[12837]<=8'd170;
		data_a[12838]<=8'd171;
		data_a[12839]<=8'd178;
		data_a[12840]<=8'd179;
		data_a[12841]<=8'd187;
		data_a[12842]<=8'd183;
		data_a[12843]<=8'd181;
		data_a[12844]<=8'd174;
		data_a[12845]<=8'd169;
		data_a[12846]<=8'd164;
		data_a[12847]<=8'd157;
		data_a[12848]<=8'd151;
		data_a[12849]<=8'd134;
		data_a[12850]<=8'd118;
		data_a[12851]<=8'd117;
		data_a[12852]<=8'd115;
		data_a[12853]<=8'd113;
		data_a[12854]<=8'd112;
		data_a[12855]<=8'd111;
		data_a[12856]<=8'd107;
		data_a[12857]<=8'd80;
		data_a[12858]<=8'd84;
		data_a[12859]<=8'd97;
		data_a[12860]<=8'd103;
		data_a[12861]<=8'd141;
		data_a[12862]<=8'd169;
		data_a[12863]<=8'd175;
		data_a[12864]<=8'd167;
		data_a[12865]<=8'd144;
		data_a[12866]<=8'd127;
		data_a[12867]<=8'd130;
		data_a[12868]<=8'd142;
		data_a[12869]<=8'd149;
		data_a[12870]<=8'd153;
		data_a[12871]<=8'd158;
		data_a[12872]<=8'd164;
		data_a[12873]<=8'd162;
		data_a[12874]<=8'd162;
		data_a[12875]<=8'd161;
		data_a[12876]<=8'd151;
		data_a[12877]<=8'd148;
		data_a[12878]<=8'd109;
		data_a[12879]<=8'd92;
		data_a[12880]<=8'd101;
		data_a[12881]<=8'd144;
		data_a[12882]<=8'd212;
		data_a[12883]<=8'd197;
		data_a[12884]<=8'd229;
		data_a[12885]<=8'd230;
		data_a[12886]<=8'd231;
		data_a[12887]<=8'd232;
		data_a[12888]<=8'd233;
		data_a[12889]<=8'd233;
		data_a[12890]<=8'd233;
		data_a[12891]<=8'd233;
		data_a[12892]<=8'd234;
		data_a[12893]<=8'd235;
		data_a[12894]<=8'd237;
		data_a[12895]<=8'd238;
		data_a[12896]<=8'd239;
		data_a[12897]<=8'd239;
		data_a[12898]<=8'd240;
		data_a[12899]<=8'd241;
		data_a[12900]<=8'd253;
		data_a[12901]<=8'd91;
		data_a[12902]<=8'd88;
		data_a[12903]<=8'd90;
		data_a[12904]<=8'd96;
		data_a[12905]<=8'd82;
		data_a[12906]<=8'd86;
		data_a[12907]<=8'd87;
		data_a[12908]<=8'd73;
		data_a[12909]<=8'd128;
		data_a[12910]<=8'd136;
		data_a[12911]<=8'd128;
		data_a[12912]<=8'd135;
		data_a[12913]<=8'd147;
		data_a[12914]<=8'd134;
		data_a[12915]<=8'd147;
		data_a[12916]<=8'd149;
		data_a[12917]<=8'd154;
		data_a[12918]<=8'd157;
		data_a[12919]<=8'd154;
		data_a[12920]<=8'd57;
		data_a[12921]<=8'd63;
		data_a[12922]<=8'd57;
		data_a[12923]<=8'd54;
		data_a[12924]<=8'd79;
		data_a[12925]<=8'd64;
		data_a[12926]<=8'd69;
		data_a[12927]<=8'd69;
		data_a[12928]<=8'd97;
		data_a[12929]<=8'd110;
		data_a[12930]<=8'd71;
		data_a[12931]<=8'd101;
		data_a[12932]<=8'd97;
		data_a[12933]<=8'd84;
		data_a[12934]<=8'd63;
		data_a[12935]<=8'd68;
		data_a[12936]<=8'd82;
		data_a[12937]<=8'd107;
		data_a[12938]<=8'd77;
		data_a[12939]<=8'd87;
		data_a[12940]<=8'd67;
		data_a[12941]<=8'd95;
		data_a[12942]<=8'd83;
		data_a[12943]<=8'd85;
		data_a[12944]<=8'd102;
		data_a[12945]<=8'd70;
		data_a[12946]<=8'd61;
		data_a[12947]<=8'd80;
		data_a[12948]<=8'd57;
		data_a[12949]<=8'd65;
		data_a[12950]<=8'd102;
		data_a[12951]<=8'd83;
		data_a[12952]<=8'd76;
		data_a[12953]<=8'd76;
		data_a[12954]<=8'd74;
		data_a[12955]<=8'd75;
		data_a[12956]<=8'd71;
		data_a[12957]<=8'd81;
		data_a[12958]<=8'd85;
		data_a[12959]<=8'd96;
		data_a[12960]<=8'd114;
		data_a[12961]<=8'd107;
		data_a[12962]<=8'd99;
		data_a[12963]<=8'd103;
		data_a[12964]<=8'd48;
		data_a[12965]<=8'd56;
		data_a[12966]<=8'd73;
		data_a[12967]<=8'd54;
		data_a[12968]<=8'd57;
		data_a[12969]<=8'd61;
		data_a[12970]<=8'd70;
		data_a[12971]<=8'd105;
		data_a[12972]<=8'd176;
		data_a[12973]<=8'd184;
		data_a[12974]<=8'd193;
		data_a[12975]<=8'd195;
		data_a[12976]<=8'd184;
		data_a[12977]<=8'd205;
		data_a[12978]<=8'd212;
		data_a[12979]<=8'd204;
		data_a[12980]<=8'd211;
		data_a[12981]<=8'd213;
		data_a[12982]<=8'd83;
		data_a[12983]<=8'd134;
		data_a[12984]<=8'd152;
		data_a[12985]<=8'd156;
		data_a[12986]<=8'd160;
		data_a[12987]<=8'd168;
		data_a[12988]<=8'd174;
		data_a[12989]<=8'd184;
		data_a[12990]<=8'd184;
		data_a[12991]<=8'd188;
		data_a[12992]<=8'd183;
		data_a[12993]<=8'd183;
		data_a[12994]<=8'd180;
		data_a[12995]<=8'd174;
		data_a[12996]<=8'd157;
		data_a[12997]<=8'd147;
		data_a[12998]<=8'd131;
		data_a[12999]<=8'd121;
		data_a[13000]<=8'd74;
		data_a[13001]<=8'd50;
		data_a[13002]<=8'd92;
		data_a[13003]<=8'd110;
		data_a[13004]<=8'd98;
		data_a[13005]<=8'd111;
		data_a[13006]<=8'd104;
		data_a[13007]<=8'd98;
		data_a[13008]<=8'd90;
		data_a[13009]<=8'd79;
		data_a[13010]<=8'd83;
		data_a[13011]<=8'd155;
		data_a[13012]<=8'd167;
		data_a[13013]<=8'd172;
		data_a[13014]<=8'd177;
		data_a[13015]<=8'd164;
		data_a[13016]<=8'd138;
		data_a[13017]<=8'd120;
		data_a[13018]<=8'd138;
		data_a[13019]<=8'd144;
		data_a[13020]<=8'd148;
		data_a[13021]<=8'd158;
		data_a[13022]<=8'd160;
		data_a[13023]<=8'd160;
		data_a[13024]<=8'd158;
		data_a[13025]<=8'd151;
		data_a[13026]<=8'd139;
		data_a[13027]<=8'd131;
		data_a[13028]<=8'd109;
		data_a[13029]<=8'd91;
		data_a[13030]<=8'd94;
		data_a[13031]<=8'd125;
		data_a[13032]<=8'd209;
		data_a[13033]<=8'd197;
		data_a[13034]<=8'd233;
		data_a[13035]<=8'd227;
		data_a[13036]<=8'd232;
		data_a[13037]<=8'd233;
		data_a[13038]<=8'd234;
		data_a[13039]<=8'd234;
		data_a[13040]<=8'd233;
		data_a[13041]<=8'd234;
		data_a[13042]<=8'd235;
		data_a[13043]<=8'd237;
		data_a[13044]<=8'd237;
		data_a[13045]<=8'd238;
		data_a[13046]<=8'd239;
		data_a[13047]<=8'd239;
		data_a[13048]<=8'd240;
		data_a[13049]<=8'd241;
		data_a[13050]<=8'd255;
		data_a[13051]<=8'd87;
		data_a[13052]<=8'd88;
		data_a[13053]<=8'd89;
		data_a[13054]<=8'd89;
		data_a[13055]<=8'd87;
		data_a[13056]<=8'd86;
		data_a[13057]<=8'd81;
		data_a[13058]<=8'd74;
		data_a[13059]<=8'd69;
		data_a[13060]<=8'd62;
		data_a[13061]<=8'd142;
		data_a[13062]<=8'd134;
		data_a[13063]<=8'd137;
		data_a[13064]<=8'd136;
		data_a[13065]<=8'd136;
		data_a[13066]<=8'd149;
		data_a[13067]<=8'd153;
		data_a[13068]<=8'd152;
		data_a[13069]<=8'd140;
		data_a[13070]<=8'd61;
		data_a[13071]<=8'd55;
		data_a[13072]<=8'd53;
		data_a[13073]<=8'd48;
		data_a[13074]<=8'd72;
		data_a[13075]<=8'd90;
		data_a[13076]<=8'd82;
		data_a[13077]<=8'd57;
		data_a[13078]<=8'd130;
		data_a[13079]<=8'd119;
		data_a[13080]<=8'd70;
		data_a[13081]<=8'd99;
		data_a[13082]<=8'd95;
		data_a[13083]<=8'd86;
		data_a[13084]<=8'd84;
		data_a[13085]<=8'd88;
		data_a[13086]<=8'd95;
		data_a[13087]<=8'd124;
		data_a[13088]<=8'd73;
		data_a[13089]<=8'd73;
		data_a[13090]<=8'd89;
		data_a[13091]<=8'd103;
		data_a[13092]<=8'd80;
		data_a[13093]<=8'd95;
		data_a[13094]<=8'd109;
		data_a[13095]<=8'd52;
		data_a[13096]<=8'd74;
		data_a[13097]<=8'd87;
		data_a[13098]<=8'd80;
		data_a[13099]<=8'd81;
		data_a[13100]<=8'd92;
		data_a[13101]<=8'd90;
		data_a[13102]<=8'd77;
		data_a[13103]<=8'd76;
		data_a[13104]<=8'd71;
		data_a[13105]<=8'd68;
		data_a[13106]<=8'd75;
		data_a[13107]<=8'd71;
		data_a[13108]<=8'd71;
		data_a[13109]<=8'd92;
		data_a[13110]<=8'd108;
		data_a[13111]<=8'd112;
		data_a[13112]<=8'd116;
		data_a[13113]<=8'd100;
		data_a[13114]<=8'd48;
		data_a[13115]<=8'd61;
		data_a[13116]<=8'd57;
		data_a[13117]<=8'd61;
		data_a[13118]<=8'd53;
		data_a[13119]<=8'd64;
		data_a[13120]<=8'd85;
		data_a[13121]<=8'd119;
		data_a[13122]<=8'd149;
		data_a[13123]<=8'd183;
		data_a[13124]<=8'd195;
		data_a[13125]<=8'd195;
		data_a[13126]<=8'd193;
		data_a[13127]<=8'd210;
		data_a[13128]<=8'd212;
		data_a[13129]<=8'd213;
		data_a[13130]<=8'd210;
		data_a[13131]<=8'd208;
		data_a[13132]<=8'd77;
		data_a[13133]<=8'd139;
		data_a[13134]<=8'd144;
		data_a[13135]<=8'd159;
		data_a[13136]<=8'd158;
		data_a[13137]<=8'd160;
		data_a[13138]<=8'd171;
		data_a[13139]<=8'd183;
		data_a[13140]<=8'd190;
		data_a[13141]<=8'd188;
		data_a[13142]<=8'd191;
		data_a[13143]<=8'd184;
		data_a[13144]<=8'd180;
		data_a[13145]<=8'd164;
		data_a[13146]<=8'd157;
		data_a[13147]<=8'd139;
		data_a[13148]<=8'd123;
		data_a[13149]<=8'd110;
		data_a[13150]<=8'd75;
		data_a[13151]<=8'd72;
		data_a[13152]<=8'd104;
		data_a[13153]<=8'd101;
		data_a[13154]<=8'd105;
		data_a[13155]<=8'd106;
		data_a[13156]<=8'd105;
		data_a[13157]<=8'd99;
		data_a[13158]<=8'd99;
		data_a[13159]<=8'd92;
		data_a[13160]<=8'd110;
		data_a[13161]<=8'd147;
		data_a[13162]<=8'd152;
		data_a[13163]<=8'd169;
		data_a[13164]<=8'd173;
		data_a[13165]<=8'd160;
		data_a[13166]<=8'd158;
		data_a[13167]<=8'd113;
		data_a[13168]<=8'd124;
		data_a[13169]<=8'd144;
		data_a[13170]<=8'd141;
		data_a[13171]<=8'd152;
		data_a[13172]<=8'd153;
		data_a[13173]<=8'd152;
		data_a[13174]<=8'd158;
		data_a[13175]<=8'd143;
		data_a[13176]<=8'd142;
		data_a[13177]<=8'd131;
		data_a[13178]<=8'd106;
		data_a[13179]<=8'd89;
		data_a[13180]<=8'd100;
		data_a[13181]<=8'd110;
		data_a[13182]<=8'd182;
		data_a[13183]<=8'd198;
		data_a[13184]<=8'd236;
		data_a[13185]<=8'd231;
		data_a[13186]<=8'd232;
		data_a[13187]<=8'd233;
		data_a[13188]<=8'd234;
		data_a[13189]<=8'd234;
		data_a[13190]<=8'd234;
		data_a[13191]<=8'd235;
		data_a[13192]<=8'd236;
		data_a[13193]<=8'd238;
		data_a[13194]<=8'd238;
		data_a[13195]<=8'd240;
		data_a[13196]<=8'd240;
		data_a[13197]<=8'd240;
		data_a[13198]<=8'd241;
		data_a[13199]<=8'd242;
		data_a[13200]<=8'd255;
		data_a[13201]<=8'd84;
		data_a[13202]<=8'd87;
		data_a[13203]<=8'd87;
		data_a[13204]<=8'd86;
		data_a[13205]<=8'd86;
		data_a[13206]<=8'd86;
		data_a[13207]<=8'd85;
		data_a[13208]<=8'd66;
		data_a[13209]<=8'd72;
		data_a[13210]<=8'd59;
		data_a[13211]<=8'd74;
		data_a[13212]<=8'd72;
		data_a[13213]<=8'd111;
		data_a[13214]<=8'd127;
		data_a[13215]<=8'd128;
		data_a[13216]<=8'd123;
		data_a[13217]<=8'd142;
		data_a[13218]<=8'd142;
		data_a[13219]<=8'd121;
		data_a[13220]<=8'd68;
		data_a[13221]<=8'd56;
		data_a[13222]<=8'd55;
		data_a[13223]<=8'd61;
		data_a[13224]<=8'd77;
		data_a[13225]<=8'd92;
		data_a[13226]<=8'd77;
		data_a[13227]<=8'd65;
		data_a[13228]<=8'd138;
		data_a[13229]<=8'd135;
		data_a[13230]<=8'd65;
		data_a[13231]<=8'd116;
		data_a[13232]<=8'd107;
		data_a[13233]<=8'd98;
		data_a[13234]<=8'd100;
		data_a[13235]<=8'd95;
		data_a[13236]<=8'd99;
		data_a[13237]<=8'd98;
		data_a[13238]<=8'd100;
		data_a[13239]<=8'd86;
		data_a[13240]<=8'd93;
		data_a[13241]<=8'd86;
		data_a[13242]<=8'd97;
		data_a[13243]<=8'd94;
		data_a[13244]<=8'd105;
		data_a[13245]<=8'd53;
		data_a[13246]<=8'd69;
		data_a[13247]<=8'd108;
		data_a[13248]<=8'd91;
		data_a[13249]<=8'd63;
		data_a[13250]<=8'd91;
		data_a[13251]<=8'd86;
		data_a[13252]<=8'd77;
		data_a[13253]<=8'd77;
		data_a[13254]<=8'd70;
		data_a[13255]<=8'd75;
		data_a[13256]<=8'd69;
		data_a[13257]<=8'd72;
		data_a[13258]<=8'd72;
		data_a[13259]<=8'd68;
		data_a[13260]<=8'd98;
		data_a[13261]<=8'd117;
		data_a[13262]<=8'd116;
		data_a[13263]<=8'd100;
		data_a[13264]<=8'd52;
		data_a[13265]<=8'd95;
		data_a[13266]<=8'd65;
		data_a[13267]<=8'd54;
		data_a[13268]<=8'd61;
		data_a[13269]<=8'd65;
		data_a[13270]<=8'd79;
		data_a[13271]<=8'd125;
		data_a[13272]<=8'd148;
		data_a[13273]<=8'd197;
		data_a[13274]<=8'd199;
		data_a[13275]<=8'd200;
		data_a[13276]<=8'd193;
		data_a[13277]<=8'd214;
		data_a[13278]<=8'd214;
		data_a[13279]<=8'd211;
		data_a[13280]<=8'd211;
		data_a[13281]<=8'd217;
		data_a[13282]<=8'd73;
		data_a[13283]<=8'd131;
		data_a[13284]<=8'd143;
		data_a[13285]<=8'd153;
		data_a[13286]<=8'd152;
		data_a[13287]<=8'd168;
		data_a[13288]<=8'd176;
		data_a[13289]<=8'd182;
		data_a[13290]<=8'd184;
		data_a[13291]<=8'd190;
		data_a[13292]<=8'd187;
		data_a[13293]<=8'd179;
		data_a[13294]<=8'd176;
		data_a[13295]<=8'd166;
		data_a[13296]<=8'd160;
		data_a[13297]<=8'd146;
		data_a[13298]<=8'd118;
		data_a[13299]<=8'd111;
		data_a[13300]<=8'd90;
		data_a[13301]<=8'd100;
		data_a[13302]<=8'd107;
		data_a[13303]<=8'd105;
		data_a[13304]<=8'd110;
		data_a[13305]<=8'd108;
		data_a[13306]<=8'd105;
		data_a[13307]<=8'd100;
		data_a[13308]<=8'd96;
		data_a[13309]<=8'd94;
		data_a[13310]<=8'd128;
		data_a[13311]<=8'd125;
		data_a[13312]<=8'd128;
		data_a[13313]<=8'd152;
		data_a[13314]<=8'd154;
		data_a[13315]<=8'd154;
		data_a[13316]<=8'd143;
		data_a[13317]<=8'd117;
		data_a[13318]<=8'd108;
		data_a[13319]<=8'd129;
		data_a[13320]<=8'd140;
		data_a[13321]<=8'd151;
		data_a[13322]<=8'd154;
		data_a[13323]<=8'd155;
		data_a[13324]<=8'd151;
		data_a[13325]<=8'd142;
		data_a[13326]<=8'd132;
		data_a[13327]<=8'd119;
		data_a[13328]<=8'd107;
		data_a[13329]<=8'd89;
		data_a[13330]<=8'd96;
		data_a[13331]<=8'd105;
		data_a[13332]<=8'd171;
		data_a[13333]<=8'd214;
		data_a[13334]<=8'd237;
		data_a[13335]<=8'd235;
		data_a[13336]<=8'd235;
		data_a[13337]<=8'd235;
		data_a[13338]<=8'd235;
		data_a[13339]<=8'd237;
		data_a[13340]<=8'd237;
		data_a[13341]<=8'd237;
		data_a[13342]<=8'd238;
		data_a[13343]<=8'd239;
		data_a[13344]<=8'd238;
		data_a[13345]<=8'd239;
		data_a[13346]<=8'd240;
		data_a[13347]<=8'd241;
		data_a[13348]<=8'd242;
		data_a[13349]<=8'd242;
		data_a[13350]<=8'd253;
		data_a[13351]<=8'd81;
		data_a[13352]<=8'd87;
		data_a[13353]<=8'd89;
		data_a[13354]<=8'd89;
		data_a[13355]<=8'd87;
		data_a[13356]<=8'd81;
		data_a[13357]<=8'd76;
		data_a[13358]<=8'd69;
		data_a[13359]<=8'd61;
		data_a[13360]<=8'd64;
		data_a[13361]<=8'd73;
		data_a[13362]<=8'd73;
		data_a[13363]<=8'd68;
		data_a[13364]<=8'd75;
		data_a[13365]<=8'd94;
		data_a[13366]<=8'd129;
		data_a[13367]<=8'd126;
		data_a[13368]<=8'd119;
		data_a[13369]<=8'd113;
		data_a[13370]<=8'd69;
		data_a[13371]<=8'd50;
		data_a[13372]<=8'd46;
		data_a[13373]<=8'd60;
		data_a[13374]<=8'd85;
		data_a[13375]<=8'd114;
		data_a[13376]<=8'd92;
		data_a[13377]<=8'd78;
		data_a[13378]<=8'd132;
		data_a[13379]<=8'd140;
		data_a[13380]<=8'd68;
		data_a[13381]<=8'd123;
		data_a[13382]<=8'd112;
		data_a[13383]<=8'd116;
		data_a[13384]<=8'd103;
		data_a[13385]<=8'd98;
		data_a[13386]<=8'd109;
		data_a[13387]<=8'd117;
		data_a[13388]<=8'd97;
		data_a[13389]<=8'd86;
		data_a[13390]<=8'd92;
		data_a[13391]<=8'd95;
		data_a[13392]<=8'd102;
		data_a[13393]<=8'd108;
		data_a[13394]<=8'd101;
		data_a[13395]<=8'd55;
		data_a[13396]<=8'd99;
		data_a[13397]<=8'd137;
		data_a[13398]<=8'd123;
		data_a[13399]<=8'd56;
		data_a[13400]<=8'd91;
		data_a[13401]<=8'd85;
		data_a[13402]<=8'd75;
		data_a[13403]<=8'd91;
		data_a[13404]<=8'd66;
		data_a[13405]<=8'd77;
		data_a[13406]<=8'd65;
		data_a[13407]<=8'd108;
		data_a[13408]<=8'd69;
		data_a[13409]<=8'd73;
		data_a[13410]<=8'd76;
		data_a[13411]<=8'd106;
		data_a[13412]<=8'd127;
		data_a[13413]<=8'd115;
		data_a[13414]<=8'd46;
		data_a[13415]<=8'd64;
		data_a[13416]<=8'd68;
		data_a[13417]<=8'd67;
		data_a[13418]<=8'd64;
		data_a[13419]<=8'd67;
		data_a[13420]<=8'd92;
		data_a[13421]<=8'd96;
		data_a[13422]<=8'd152;
		data_a[13423]<=8'd199;
		data_a[13424]<=8'd201;
		data_a[13425]<=8'd205;
		data_a[13426]<=8'd201;
		data_a[13427]<=8'd217;
		data_a[13428]<=8'd214;
		data_a[13429]<=8'd214;
		data_a[13430]<=8'd218;
		data_a[13431]<=8'd215;
		data_a[13432]<=8'd95;
		data_a[13433]<=8'd120;
		data_a[13434]<=8'd140;
		data_a[13435]<=8'd155;
		data_a[13436]<=8'd153;
		data_a[13437]<=8'd165;
		data_a[13438]<=8'd173;
		data_a[13439]<=8'd184;
		data_a[13440]<=8'd188;
		data_a[13441]<=8'd186;
		data_a[13442]<=8'd182;
		data_a[13443]<=8'd182;
		data_a[13444]<=8'd179;
		data_a[13445]<=8'd168;
		data_a[13446]<=8'd157;
		data_a[13447]<=8'd151;
		data_a[13448]<=8'd121;
		data_a[13449]<=8'd106;
		data_a[13450]<=8'd93;
		data_a[13451]<=8'd94;
		data_a[13452]<=8'd100;
		data_a[13453]<=8'd107;
		data_a[13454]<=8'd115;
		data_a[13455]<=8'd112;
		data_a[13456]<=8'd105;
		data_a[13457]<=8'd93;
		data_a[13458]<=8'd95;
		data_a[13459]<=8'd96;
		data_a[13460]<=8'd104;
		data_a[13461]<=8'd110;
		data_a[13462]<=8'd139;
		data_a[13463]<=8'd139;
		data_a[13464]<=8'd138;
		data_a[13465]<=8'd121;
		data_a[13466]<=8'd124;
		data_a[13467]<=8'd119;
		data_a[13468]<=8'd87;
		data_a[13469]<=8'd116;
		data_a[13470]<=8'd134;
		data_a[13471]<=8'd141;
		data_a[13472]<=8'd151;
		data_a[13473]<=8'd154;
		data_a[13474]<=8'd150;
		data_a[13475]<=8'd127;
		data_a[13476]<=8'd124;
		data_a[13477]<=8'd114;
		data_a[13478]<=8'd97;
		data_a[13479]<=8'd87;
		data_a[13480]<=8'd92;
		data_a[13481]<=8'd100;
		data_a[13482]<=8'd180;
		data_a[13483]<=8'd215;
		data_a[13484]<=8'd235;
		data_a[13485]<=8'd231;
		data_a[13486]<=8'd235;
		data_a[13487]<=8'd235;
		data_a[13488]<=8'd235;
		data_a[13489]<=8'd237;
		data_a[13490]<=8'd238;
		data_a[13491]<=8'd238;
		data_a[13492]<=8'd238;
		data_a[13493]<=8'd239;
		data_a[13494]<=8'd241;
		data_a[13495]<=8'd241;
		data_a[13496]<=8'd242;
		data_a[13497]<=8'd243;
		data_a[13498]<=8'd244;
		data_a[13499]<=8'd243;
		data_a[13500]<=8'd255;
		data_a[13501]<=8'd78;
		data_a[13502]<=8'd79;
		data_a[13503]<=8'd79;
		data_a[13504]<=8'd82;
		data_a[13505]<=8'd86;
		data_a[13506]<=8'd86;
		data_a[13507]<=8'd84;
		data_a[13508]<=8'd68;
		data_a[13509]<=8'd65;
		data_a[13510]<=8'd66;
		data_a[13511]<=8'd76;
		data_a[13512]<=8'd73;
		data_a[13513]<=8'd65;
		data_a[13514]<=8'd53;
		data_a[13515]<=8'd74;
		data_a[13516]<=8'd65;
		data_a[13517]<=8'd87;
		data_a[13518]<=8'd115;
		data_a[13519]<=8'd115;
		data_a[13520]<=8'd63;
		data_a[13521]<=8'd52;
		data_a[13522]<=8'd54;
		data_a[13523]<=8'd51;
		data_a[13524]<=8'd82;
		data_a[13525]<=8'd107;
		data_a[13526]<=8'd90;
		data_a[13527]<=8'd84;
		data_a[13528]<=8'd136;
		data_a[13529]<=8'd144;
		data_a[13530]<=8'd55;
		data_a[13531]<=8'd135;
		data_a[13532]<=8'd128;
		data_a[13533]<=8'd116;
		data_a[13534]<=8'd116;
		data_a[13535]<=8'd106;
		data_a[13536]<=8'd104;
		data_a[13537]<=8'd103;
		data_a[13538]<=8'd104;
		data_a[13539]<=8'd102;
		data_a[13540]<=8'd102;
		data_a[13541]<=8'd101;
		data_a[13542]<=8'd108;
		data_a[13543]<=8'd114;
		data_a[13544]<=8'd80;
		data_a[13545]<=8'd58;
		data_a[13546]<=8'd133;
		data_a[13547]<=8'd157;
		data_a[13548]<=8'd140;
		data_a[13549]<=8'd77;
		data_a[13550]<=8'd64;
		data_a[13551]<=8'd90;
		data_a[13552]<=8'd78;
		data_a[13553]<=8'd81;
		data_a[13554]<=8'd94;
		data_a[13555]<=8'd68;
		data_a[13556]<=8'd67;
		data_a[13557]<=8'd128;
		data_a[13558]<=8'd62;
		data_a[13559]<=8'd59;
		data_a[13560]<=8'd78;
		data_a[13561]<=8'd107;
		data_a[13562]<=8'd122;
		data_a[13563]<=8'd128;
		data_a[13564]<=8'd53;
		data_a[13565]<=8'd67;
		data_a[13566]<=8'd73;
		data_a[13567]<=8'd63;
		data_a[13568]<=8'd69;
		data_a[13569]<=8'd76;
		data_a[13570]<=8'd98;
		data_a[13571]<=8'd108;
		data_a[13572]<=8'd165;
		data_a[13573]<=8'd202;
		data_a[13574]<=8'd202;
		data_a[13575]<=8'd208;
		data_a[13576]<=8'd206;
		data_a[13577]<=8'd218;
		data_a[13578]<=8'd215;
		data_a[13579]<=8'd218;
		data_a[13580]<=8'd214;
		data_a[13581]<=8'd216;
		data_a[13582]<=8'd100;
		data_a[13583]<=8'd115;
		data_a[13584]<=8'd139;
		data_a[13585]<=8'd145;
		data_a[13586]<=8'd156;
		data_a[13587]<=8'd164;
		data_a[13588]<=8'd169;
		data_a[13589]<=8'd178;
		data_a[13590]<=8'd186;
		data_a[13591]<=8'd184;
		data_a[13592]<=8'd182;
		data_a[13593]<=8'd182;
		data_a[13594]<=8'd174;
		data_a[13595]<=8'd164;
		data_a[13596]<=8'd166;
		data_a[13597]<=8'd160;
		data_a[13598]<=8'd140;
		data_a[13599]<=8'd95;
		data_a[13600]<=8'd74;
		data_a[13601]<=8'd92;
		data_a[13602]<=8'd97;
		data_a[13603]<=8'd102;
		data_a[13604]<=8'd103;
		data_a[13605]<=8'd111;
		data_a[13606]<=8'd99;
		data_a[13607]<=8'd95;
		data_a[13608]<=8'd89;
		data_a[13609]<=8'd86;
		data_a[13610]<=8'd88;
		data_a[13611]<=8'd91;
		data_a[13612]<=8'd115;
		data_a[13613]<=8'd121;
		data_a[13614]<=8'd119;
		data_a[13615]<=8'd106;
		data_a[13616]<=8'd100;
		data_a[13617]<=8'd96;
		data_a[13618]<=8'd85;
		data_a[13619]<=8'd108;
		data_a[13620]<=8'd130;
		data_a[13621]<=8'd144;
		data_a[13622]<=8'd139;
		data_a[13623]<=8'd143;
		data_a[13624]<=8'd148;
		data_a[13625]<=8'd124;
		data_a[13626]<=8'd109;
		data_a[13627]<=8'd107;
		data_a[13628]<=8'd97;
		data_a[13629]<=8'd92;
		data_a[13630]<=8'd84;
		data_a[13631]<=8'd106;
		data_a[13632]<=8'd144;
		data_a[13633]<=8'd198;
		data_a[13634]<=8'd237;
		data_a[13635]<=8'd234;
		data_a[13636]<=8'd236;
		data_a[13637]<=8'd235;
		data_a[13638]<=8'd236;
		data_a[13639]<=8'd237;
		data_a[13640]<=8'd238;
		data_a[13641]<=8'd238;
		data_a[13642]<=8'd239;
		data_a[13643]<=8'd240;
		data_a[13644]<=8'd242;
		data_a[13645]<=8'd243;
		data_a[13646]<=8'd243;
		data_a[13647]<=8'd244;
		data_a[13648]<=8'd245;
		data_a[13649]<=8'd244;
		data_a[13650]<=8'd255;
		data_a[13651]<=8'd79;
		data_a[13652]<=8'd78;
		data_a[13653]<=8'd77;
		data_a[13654]<=8'd79;
		data_a[13655]<=8'd82;
		data_a[13656]<=8'd81;
		data_a[13657]<=8'd78;
		data_a[13658]<=8'd69;
		data_a[13659]<=8'd62;
		data_a[13660]<=8'd60;
		data_a[13661]<=8'd63;
		data_a[13662]<=8'd82;
		data_a[13663]<=8'd82;
		data_a[13664]<=8'd70;
		data_a[13665]<=8'd65;
		data_a[13666]<=8'd67;
		data_a[13667]<=8'd59;
		data_a[13668]<=8'd56;
		data_a[13669]<=8'd73;
		data_a[13670]<=8'd66;
		data_a[13671]<=8'd55;
		data_a[13672]<=8'd43;
		data_a[13673]<=8'd51;
		data_a[13674]<=8'd86;
		data_a[13675]<=8'd100;
		data_a[13676]<=8'd90;
		data_a[13677]<=8'd87;
		data_a[13678]<=8'd143;
		data_a[13679]<=8'd140;
		data_a[13680]<=8'd63;
		data_a[13681]<=8'd147;
		data_a[13682]<=8'd135;
		data_a[13683]<=8'd129;
		data_a[13684]<=8'd130;
		data_a[13685]<=8'd113;
		data_a[13686]<=8'd116;
		data_a[13687]<=8'd107;
		data_a[13688]<=8'd104;
		data_a[13689]<=8'd106;
		data_a[13690]<=8'd103;
		data_a[13691]<=8'd113;
		data_a[13692]<=8'd126;
		data_a[13693]<=8'd114;
		data_a[13694]<=8'd77;
		data_a[13695]<=8'd86;
		data_a[13696]<=8'd160;
		data_a[13697]<=8'd199;
		data_a[13698]<=8'd161;
		data_a[13699]<=8'd128;
		data_a[13700]<=8'd40;
		data_a[13701]<=8'd95;
		data_a[13702]<=8'd81;
		data_a[13703]<=8'd87;
		data_a[13704]<=8'd87;
		data_a[13705]<=8'd82;
		data_a[13706]<=8'd78;
		data_a[13707]<=8'd64;
		data_a[13708]<=8'd70;
		data_a[13709]<=8'd68;
		data_a[13710]<=8'd67;
		data_a[13711]<=8'd89;
		data_a[13712]<=8'd122;
		data_a[13713]<=8'd140;
		data_a[13714]<=8'd67;
		data_a[13715]<=8'd74;
		data_a[13716]<=8'd65;
		data_a[13717]<=8'd73;
		data_a[13718]<=8'd78;
		data_a[13719]<=8'd80;
		data_a[13720]<=8'd140;
		data_a[13721]<=8'd102;
		data_a[13722]<=8'd188;
		data_a[13723]<=8'd207;
		data_a[13724]<=8'd204;
		data_a[13725]<=8'd209;
		data_a[13726]<=8'd204;
		data_a[13727]<=8'd218;
		data_a[13728]<=8'd219;
		data_a[13729]<=8'd222;
		data_a[13730]<=8'd220;
		data_a[13731]<=8'd219;
		data_a[13732]<=8'd113;
		data_a[13733]<=8'd97;
		data_a[13734]<=8'd129;
		data_a[13735]<=8'd153;
		data_a[13736]<=8'd149;
		data_a[13737]<=8'd160;
		data_a[13738]<=8'd171;
		data_a[13739]<=8'd171;
		data_a[13740]<=8'd179;
		data_a[13741]<=8'd182;
		data_a[13742]<=8'd184;
		data_a[13743]<=8'd179;
		data_a[13744]<=8'd166;
		data_a[13745]<=8'd163;
		data_a[13746]<=8'd164;
		data_a[13747]<=8'd179;
		data_a[13748]<=8'd152;
		data_a[13749]<=8'd125;
		data_a[13750]<=8'd103;
		data_a[13751]<=8'd89;
		data_a[13752]<=8'd86;
		data_a[13753]<=8'd88;
		data_a[13754]<=8'd104;
		data_a[13755]<=8'd98;
		data_a[13756]<=8'd91;
		data_a[13757]<=8'd90;
		data_a[13758]<=8'd82;
		data_a[13759]<=8'd93;
		data_a[13760]<=8'd83;
		data_a[13761]<=8'd80;
		data_a[13762]<=8'd93;
		data_a[13763]<=8'd103;
		data_a[13764]<=8'd103;
		data_a[13765]<=8'd109;
		data_a[13766]<=8'd96;
		data_a[13767]<=8'd91;
		data_a[13768]<=8'd100;
		data_a[13769]<=8'd96;
		data_a[13770]<=8'd115;
		data_a[13771]<=8'd136;
		data_a[13772]<=8'd146;
		data_a[13773]<=8'd143;
		data_a[13774]<=8'd135;
		data_a[13775]<=8'd112;
		data_a[13776]<=8'd107;
		data_a[13777]<=8'd100;
		data_a[13778]<=8'd84;
		data_a[13779]<=8'd92;
		data_a[13780]<=8'd75;
		data_a[13781]<=8'd90;
		data_a[13782]<=8'd137;
		data_a[13783]<=8'd193;
		data_a[13784]<=8'd237;
		data_a[13785]<=8'd233;
		data_a[13786]<=8'd237;
		data_a[13787]<=8'd236;
		data_a[13788]<=8'd237;
		data_a[13789]<=8'd238;
		data_a[13790]<=8'd239;
		data_a[13791]<=8'd239;
		data_a[13792]<=8'd239;
		data_a[13793]<=8'd240;
		data_a[13794]<=8'd241;
		data_a[13795]<=8'd242;
		data_a[13796]<=8'd243;
		data_a[13797]<=8'd244;
		data_a[13798]<=8'd245;
		data_a[13799]<=8'd245;
		data_a[13800]<=8'd253;
		data_a[13801]<=8'd76;
		data_a[13802]<=8'd76;
		data_a[13803]<=8'd76;
		data_a[13804]<=8'd76;
		data_a[13805]<=8'd77;
		data_a[13806]<=8'd74;
		data_a[13807]<=8'd71;
		data_a[13808]<=8'd61;
		data_a[13809]<=8'd63;
		data_a[13810]<=8'd61;
		data_a[13811]<=8'd78;
		data_a[13812]<=8'd69;
		data_a[13813]<=8'd70;
		data_a[13814]<=8'd70;
		data_a[13815]<=8'd76;
		data_a[13816]<=8'd69;
		data_a[13817]<=8'd66;
		data_a[13818]<=8'd62;
		data_a[13819]<=8'd67;
		data_a[13820]<=8'd61;
		data_a[13821]<=8'd63;
		data_a[13822]<=8'd54;
		data_a[13823]<=8'd43;
		data_a[13824]<=8'd111;
		data_a[13825]<=8'd106;
		data_a[13826]<=8'd87;
		data_a[13827]<=8'd82;
		data_a[13828]<=8'd145;
		data_a[13829]<=8'd144;
		data_a[13830]<=8'd127;
		data_a[13831]<=8'd165;
		data_a[13832]<=8'd148;
		data_a[13833]<=8'd148;
		data_a[13834]<=8'd143;
		data_a[13835]<=8'd131;
		data_a[13836]<=8'd120;
		data_a[13837]<=8'd124;
		data_a[13838]<=8'd120;
		data_a[13839]<=8'd120;
		data_a[13840]<=8'd128;
		data_a[13841]<=8'd131;
		data_a[13842]<=8'd130;
		data_a[13843]<=8'd112;
		data_a[13844]<=8'd58;
		data_a[13845]<=8'd143;
		data_a[13846]<=8'd173;
		data_a[13847]<=8'd190;
		data_a[13848]<=8'd171;
		data_a[13849]<=8'd135;
		data_a[13850]<=8'd58;
		data_a[13851]<=8'd99;
		data_a[13852]<=8'd96;
		data_a[13853]<=8'd83;
		data_a[13854]<=8'd90;
		data_a[13855]<=8'd82;
		data_a[13856]<=8'd84;
		data_a[13857]<=8'd87;
		data_a[13858]<=8'd90;
		data_a[13859]<=8'd81;
		data_a[13860]<=8'd88;
		data_a[13861]<=8'd89;
		data_a[13862]<=8'd133;
		data_a[13863]<=8'd136;
		data_a[13864]<=8'd116;
		data_a[13865]<=8'd87;
		data_a[13866]<=8'd77;
		data_a[13867]<=8'd69;
		data_a[13868]<=8'd71;
		data_a[13869]<=8'd87;
		data_a[13870]<=8'd155;
		data_a[13871]<=8'd97;
		data_a[13872]<=8'd207;
		data_a[13873]<=8'd209;
		data_a[13874]<=8'd206;
		data_a[13875]<=8'd213;
		data_a[13876]<=8'd204;
		data_a[13877]<=8'd219;
		data_a[13878]<=8'd224;
		data_a[13879]<=8'd223;
		data_a[13880]<=8'd222;
		data_a[13881]<=8'd216;
		data_a[13882]<=8'd121;
		data_a[13883]<=8'd79;
		data_a[13884]<=8'd131;
		data_a[13885]<=8'd139;
		data_a[13886]<=8'd147;
		data_a[13887]<=8'd167;
		data_a[13888]<=8'd172;
		data_a[13889]<=8'd170;
		data_a[13890]<=8'd176;
		data_a[13891]<=8'd179;
		data_a[13892]<=8'd180;
		data_a[13893]<=8'd174;
		data_a[13894]<=8'd166;
		data_a[13895]<=8'd172;
		data_a[13896]<=8'd175;
		data_a[13897]<=8'd171;
		data_a[13898]<=8'd153;
		data_a[13899]<=8'd134;
		data_a[13900]<=8'd93;
		data_a[13901]<=8'd83;
		data_a[13902]<=8'd81;
		data_a[13903]<=8'd80;
		data_a[13904]<=8'd88;
		data_a[13905]<=8'd95;
		data_a[13906]<=8'd71;
		data_a[13907]<=8'd78;
		data_a[13908]<=8'd71;
		data_a[13909]<=8'd72;
		data_a[13910]<=8'd79;
		data_a[13911]<=8'd71;
		data_a[13912]<=8'd87;
		data_a[13913]<=8'd87;
		data_a[13914]<=8'd98;
		data_a[13915]<=8'd100;
		data_a[13916]<=8'd89;
		data_a[13917]<=8'd94;
		data_a[13918]<=8'd91;
		data_a[13919]<=8'd87;
		data_a[13920]<=8'd89;
		data_a[13921]<=8'd127;
		data_a[13922]<=8'd149;
		data_a[13923]<=8'd139;
		data_a[13924]<=8'd139;
		data_a[13925]<=8'd107;
		data_a[13926]<=8'd97;
		data_a[13927]<=8'd99;
		data_a[13928]<=8'd85;
		data_a[13929]<=8'd92;
		data_a[13930]<=8'd83;
		data_a[13931]<=8'd90;
		data_a[13932]<=8'd134;
		data_a[13933]<=8'd213;
		data_a[13934]<=8'd238;
		data_a[13935]<=8'd236;
		data_a[13936]<=8'd238;
		data_a[13937]<=8'd237;
		data_a[13938]<=8'd238;
		data_a[13939]<=8'd239;
		data_a[13940]<=8'd240;
		data_a[13941]<=8'd239;
		data_a[13942]<=8'd240;
		data_a[13943]<=8'd241;
		data_a[13944]<=8'd241;
		data_a[13945]<=8'd242;
		data_a[13946]<=8'd243;
		data_a[13947]<=8'd244;
		data_a[13948]<=8'd245;
		data_a[13949]<=8'd245;
		data_a[13950]<=8'd254;
		data_a[13951]<=8'd76;
		data_a[13952]<=8'd74;
		data_a[13953]<=8'd71;
		data_a[13954]<=8'd71;
		data_a[13955]<=8'd74;
		data_a[13956]<=8'd75;
		data_a[13957]<=8'd74;
		data_a[13958]<=8'd70;
		data_a[13959]<=8'd55;
		data_a[13960]<=8'd61;
		data_a[13961]<=8'd71;
		data_a[13962]<=8'd79;
		data_a[13963]<=8'd63;
		data_a[13964]<=8'd74;
		data_a[13965]<=8'd65;
		data_a[13966]<=8'd61;
		data_a[13967]<=8'd70;
		data_a[13968]<=8'd59;
		data_a[13969]<=8'd58;
		data_a[13970]<=8'd68;
		data_a[13971]<=8'd66;
		data_a[13972]<=8'd48;
		data_a[13973]<=8'd48;
		data_a[13974]<=8'd105;
		data_a[13975]<=8'd104;
		data_a[13976]<=8'd83;
		data_a[13977]<=8'd90;
		data_a[13978]<=8'd140;
		data_a[13979]<=8'd138;
		data_a[13980]<=8'd153;
		data_a[13981]<=8'd63;
		data_a[13982]<=8'd170;
		data_a[13983]<=8'd154;
		data_a[13984]<=8'd156;
		data_a[13985]<=8'd157;
		data_a[13986]<=8'd142;
		data_a[13987]<=8'd130;
		data_a[13988]<=8'd135;
		data_a[13989]<=8'd134;
		data_a[13990]<=8'd137;
		data_a[13991]<=8'd129;
		data_a[13992]<=8'd131;
		data_a[13993]<=8'd99;
		data_a[13994]<=8'd67;
		data_a[13995]<=8'd154;
		data_a[13996]<=8'd176;
		data_a[13997]<=8'd195;
		data_a[13998]<=8'd182;
		data_a[13999]<=8'd145;
		data_a[14000]<=8'd40;
		data_a[14001]<=8'd106;
		data_a[14002]<=8'd107;
		data_a[14003]<=8'd100;
		data_a[14004]<=8'd73;
		data_a[14005]<=8'd76;
		data_a[14006]<=8'd79;
		data_a[14007]<=8'd78;
		data_a[14008]<=8'd86;
		data_a[14009]<=8'd95;
		data_a[14010]<=8'd114;
		data_a[14011]<=8'd116;
		data_a[14012]<=8'd122;
		data_a[14013]<=8'd127;
		data_a[14014]<=8'd144;
		data_a[14015]<=8'd67;
		data_a[14016]<=8'd73;
		data_a[14017]<=8'd91;
		data_a[14018]<=8'd77;
		data_a[14019]<=8'd89;
		data_a[14020]<=8'd136;
		data_a[14021]<=8'd162;
		data_a[14022]<=8'd211;
		data_a[14023]<=8'd208;
		data_a[14024]<=8'd209;
		data_a[14025]<=8'd216;
		data_a[14026]<=8'd208;
		data_a[14027]<=8'd222;
		data_a[14028]<=8'd226;
		data_a[14029]<=8'd221;
		data_a[14030]<=8'd221;
		data_a[14031]<=8'd227;
		data_a[14032]<=8'd109;
		data_a[14033]<=8'd84;
		data_a[14034]<=8'd128;
		data_a[14035]<=8'd147;
		data_a[14036]<=8'd148;
		data_a[14037]<=8'd158;
		data_a[14038]<=8'd162;
		data_a[14039]<=8'd171;
		data_a[14040]<=8'd177;
		data_a[14041]<=8'd177;
		data_a[14042]<=8'd175;
		data_a[14043]<=8'd170;
		data_a[14044]<=8'd168;
		data_a[14045]<=8'd177;
		data_a[14046]<=8'd174;
		data_a[14047]<=8'd185;
		data_a[14048]<=8'd143;
		data_a[14049]<=8'd129;
		data_a[14050]<=8'd97;
		data_a[14051]<=8'd80;
		data_a[14052]<=8'd82;
		data_a[14053]<=8'd76;
		data_a[14054]<=8'd74;
		data_a[14055]<=8'd92;
		data_a[14056]<=8'd80;
		data_a[14057]<=8'd74;
		data_a[14058]<=8'd74;
		data_a[14059]<=8'd70;
		data_a[14060]<=8'd70;
		data_a[14061]<=8'd80;
		data_a[14062]<=8'd78;
		data_a[14063]<=8'd84;
		data_a[14064]<=8'd88;
		data_a[14065]<=8'd82;
		data_a[14066]<=8'd77;
		data_a[14067]<=8'd81;
		data_a[14068]<=8'd76;
		data_a[14069]<=8'd86;
		data_a[14070]<=8'd82;
		data_a[14071]<=8'd108;
		data_a[14072]<=8'd141;
		data_a[14073]<=8'd151;
		data_a[14074]<=8'd129;
		data_a[14075]<=8'd111;
		data_a[14076]<=8'd99;
		data_a[14077]<=8'd101;
		data_a[14078]<=8'd88;
		data_a[14079]<=8'd82;
		data_a[14080]<=8'd84;
		data_a[14081]<=8'd87;
		data_a[14082]<=8'd116;
		data_a[14083]<=8'd224;
		data_a[14084]<=8'd231;
		data_a[14085]<=8'd235;
		data_a[14086]<=8'd238;
		data_a[14087]<=8'd238;
		data_a[14088]<=8'd238;
		data_a[14089]<=8'd240;
		data_a[14090]<=8'd240;
		data_a[14091]<=8'd240;
		data_a[14092]<=8'd241;
		data_a[14093]<=8'd242;
		data_a[14094]<=8'd243;
		data_a[14095]<=8'd243;
		data_a[14096]<=8'd244;
		data_a[14097]<=8'd245;
		data_a[14098]<=8'd245;
		data_a[14099]<=8'd245;
		data_a[14100]<=8'd255;
		data_a[14101]<=8'd80;
		data_a[14102]<=8'd80;
		data_a[14103]<=8'd77;
		data_a[14104]<=8'd76;
		data_a[14105]<=8'd75;
		data_a[14106]<=8'd72;
		data_a[14107]<=8'd67;
		data_a[14108]<=8'd64;
		data_a[14109]<=8'd56;
		data_a[14110]<=8'd60;
		data_a[14111]<=8'd70;
		data_a[14112]<=8'd68;
		data_a[14113]<=8'd69;
		data_a[14114]<=8'd70;
		data_a[14115]<=8'd63;
		data_a[14116]<=8'd71;
		data_a[14117]<=8'd66;
		data_a[14118]<=8'd55;
		data_a[14119]<=8'd57;
		data_a[14120]<=8'd64;
		data_a[14121]<=8'd71;
		data_a[14122]<=8'd61;
		data_a[14123]<=8'd52;
		data_a[14124]<=8'd105;
		data_a[14125]<=8'd94;
		data_a[14126]<=8'd95;
		data_a[14127]<=8'd83;
		data_a[14128]<=8'd143;
		data_a[14129]<=8'd144;
		data_a[14130]<=8'd141;
		data_a[14131]<=8'd152;
		data_a[14132]<=8'd45;
		data_a[14133]<=8'd130;
		data_a[14134]<=8'd181;
		data_a[14135]<=8'd166;
		data_a[14136]<=8'd160;
		data_a[14137]<=8'd146;
		data_a[14138]<=8'd150;
		data_a[14139]<=8'd144;
		data_a[14140]<=8'd129;
		data_a[14141]<=8'd134;
		data_a[14142]<=8'd123;
		data_a[14143]<=8'd65;
		data_a[14144]<=8'd125;
		data_a[14145]<=8'd165;
		data_a[14146]<=8'd183;
		data_a[14147]<=8'd184;
		data_a[14148]<=8'd187;
		data_a[14149]<=8'd155;
		data_a[14150]<=8'd115;
		data_a[14151]<=8'd64;
		data_a[14152]<=8'd99;
		data_a[14153]<=8'd90;
		data_a[14154]<=8'd101;
		data_a[14155]<=8'd78;
		data_a[14156]<=8'd79;
		data_a[14157]<=8'd90;
		data_a[14158]<=8'd99;
		data_a[14159]<=8'd115;
		data_a[14160]<=8'd117;
		data_a[14161]<=8'd123;
		data_a[14162]<=8'd126;
		data_a[14163]<=8'd82;
		data_a[14164]<=8'd137;
		data_a[14165]<=8'd109;
		data_a[14166]<=8'd69;
		data_a[14167]<=8'd78;
		data_a[14168]<=8'd84;
		data_a[14169]<=8'd91;
		data_a[14170]<=8'd141;
		data_a[14171]<=8'd210;
		data_a[14172]<=8'd210;
		data_a[14173]<=8'd211;
		data_a[14174]<=8'd212;
		data_a[14175]<=8'd217;
		data_a[14176]<=8'd213;
		data_a[14177]<=8'd225;
		data_a[14178]<=8'd225;
		data_a[14179]<=8'd223;
		data_a[14180]<=8'd218;
		data_a[14181]<=8'd232;
		data_a[14182]<=8'd138;
		data_a[14183]<=8'd79;
		data_a[14184]<=8'd112;
		data_a[14185]<=8'd137;
		data_a[14186]<=8'd146;
		data_a[14187]<=8'd152;
		data_a[14188]<=8'd153;
		data_a[14189]<=8'd169;
		data_a[14190]<=8'd175;
		data_a[14191]<=8'd174;
		data_a[14192]<=8'd172;
		data_a[14193]<=8'd167;
		data_a[14194]<=8'd168;
		data_a[14195]<=8'd174;
		data_a[14196]<=8'd178;
		data_a[14197]<=8'd165;
		data_a[14198]<=8'd131;
		data_a[14199]<=8'd113;
		data_a[14200]<=8'd86;
		data_a[14201]<=8'd74;
		data_a[14202]<=8'd71;
		data_a[14203]<=8'd74;
		data_a[14204]<=8'd66;
		data_a[14205]<=8'd84;
		data_a[14206]<=8'd71;
		data_a[14207]<=8'd68;
		data_a[14208]<=8'd83;
		data_a[14209]<=8'd72;
		data_a[14210]<=8'd70;
		data_a[14211]<=8'd69;
		data_a[14212]<=8'd75;
		data_a[14213]<=8'd85;
		data_a[14214]<=8'd75;
		data_a[14215]<=8'd74;
		data_a[14216]<=8'd75;
		data_a[14217]<=8'd75;
		data_a[14218]<=8'd76;
		data_a[14219]<=8'd82;
		data_a[14220]<=8'd75;
		data_a[14221]<=8'd101;
		data_a[14222]<=8'd139;
		data_a[14223]<=8'd150;
		data_a[14224]<=8'd121;
		data_a[14225]<=8'd106;
		data_a[14226]<=8'd90;
		data_a[14227]<=8'd108;
		data_a[14228]<=8'd82;
		data_a[14229]<=8'd85;
		data_a[14230]<=8'd82;
		data_a[14231]<=8'd80;
		data_a[14232]<=8'd140;
		data_a[14233]<=8'd234;
		data_a[14234]<=8'd235;
		data_a[14235]<=8'd240;
		data_a[14236]<=8'd239;
		data_a[14237]<=8'd238;
		data_a[14238]<=8'd239;
		data_a[14239]<=8'd240;
		data_a[14240]<=8'd241;
		data_a[14241]<=8'd241;
		data_a[14242]<=8'd241;
		data_a[14243]<=8'd242;
		data_a[14244]<=8'd244;
		data_a[14245]<=8'd244;
		data_a[14246]<=8'd245;
		data_a[14247]<=8'd246;
		data_a[14248]<=8'd246;
		data_a[14249]<=8'd246;
		data_a[14250]<=8'd254;
		data_a[14251]<=8'd79;
		data_a[14252]<=8'd80;
		data_a[14253]<=8'd79;
		data_a[14254]<=8'd79;
		data_a[14255]<=8'd78;
		data_a[14256]<=8'd75;
		data_a[14257]<=8'd70;
		data_a[14258]<=8'd62;
		data_a[14259]<=8'd59;
		data_a[14260]<=8'd64;
		data_a[14261]<=8'd69;
		data_a[14262]<=8'd63;
		data_a[14263]<=8'd72;
		data_a[14264]<=8'd69;
		data_a[14265]<=8'd70;
		data_a[14266]<=8'd65;
		data_a[14267]<=8'd66;
		data_a[14268]<=8'd58;
		data_a[14269]<=8'd55;
		data_a[14270]<=8'd60;
		data_a[14271]<=8'd69;
		data_a[14272]<=8'd66;
		data_a[14273]<=8'd62;
		data_a[14274]<=8'd121;
		data_a[14275]<=8'd98;
		data_a[14276]<=8'd86;
		data_a[14277]<=8'd87;
		data_a[14278]<=8'd140;
		data_a[14279]<=8'd147;
		data_a[14280]<=8'd148;
		data_a[14281]<=8'd160;
		data_a[14282]<=8'd171;
		data_a[14283]<=8'd134;
		data_a[14284]<=8'd68;
		data_a[14285]<=8'd57;
		data_a[14286]<=8'd92;
		data_a[14287]<=8'd117;
		data_a[14288]<=8'd126;
		data_a[14289]<=8'd121;
		data_a[14290]<=8'd113;
		data_a[14291]<=8'd87;
		data_a[14292]<=8'd62;
		data_a[14293]<=8'd97;
		data_a[14294]<=8'd159;
		data_a[14295]<=8'd172;
		data_a[14296]<=8'd179;
		data_a[14297]<=8'd191;
		data_a[14298]<=8'd182;
		data_a[14299]<=8'd160;
		data_a[14300]<=8'd130;
		data_a[14301]<=8'd56;
		data_a[14302]<=8'd107;
		data_a[14303]<=8'd98;
		data_a[14304]<=8'd104;
		data_a[14305]<=8'd96;
		data_a[14306]<=8'd99;
		data_a[14307]<=8'd106;
		data_a[14308]<=8'd116;
		data_a[14309]<=8'd126;
		data_a[14310]<=8'd118;
		data_a[14311]<=8'd122;
		data_a[14312]<=8'd138;
		data_a[14313]<=8'd48;
		data_a[14314]<=8'd146;
		data_a[14315]<=8'd116;
		data_a[14316]<=8'd79;
		data_a[14317]<=8'd85;
		data_a[14318]<=8'd111;
		data_a[14319]<=8'd106;
		data_a[14320]<=8'd171;
		data_a[14321]<=8'd208;
		data_a[14322]<=8'd211;
		data_a[14323]<=8'd218;
		data_a[14324]<=8'd216;
		data_a[14325]<=8'd216;
		data_a[14326]<=8'd217;
		data_a[14327]<=8'd228;
		data_a[14328]<=8'd226;
		data_a[14329]<=8'd228;
		data_a[14330]<=8'd226;
		data_a[14331]<=8'd224;
		data_a[14332]<=8'd89;
		data_a[14333]<=8'd82;
		data_a[14334]<=8'd96;
		data_a[14335]<=8'd136;
		data_a[14336]<=8'd137;
		data_a[14337]<=8'd149;
		data_a[14338]<=8'd155;
		data_a[14339]<=8'd168;
		data_a[14340]<=8'd168;
		data_a[14341]<=8'd169;
		data_a[14342]<=8'd170;
		data_a[14343]<=8'd165;
		data_a[14344]<=8'd168;
		data_a[14345]<=8'd174;
		data_a[14346]<=8'd167;
		data_a[14347]<=8'd166;
		data_a[14348]<=8'd125;
		data_a[14349]<=8'd93;
		data_a[14350]<=8'd83;
		data_a[14351]<=8'd77;
		data_a[14352]<=8'd71;
		data_a[14353]<=8'd70;
		data_a[14354]<=8'd69;
		data_a[14355]<=8'd72;
		data_a[14356]<=8'd74;
		data_a[14357]<=8'd63;
		data_a[14358]<=8'd76;
		data_a[14359]<=8'd73;
		data_a[14360]<=8'd70;
		data_a[14361]<=8'd67;
		data_a[14362]<=8'd73;
		data_a[14363]<=8'd79;
		data_a[14364]<=8'd78;
		data_a[14365]<=8'd77;
		data_a[14366]<=8'd69;
		data_a[14367]<=8'd69;
		data_a[14368]<=8'd72;
		data_a[14369]<=8'd75;
		data_a[14370]<=8'd76;
		data_a[14371]<=8'd84;
		data_a[14372]<=8'd140;
		data_a[14373]<=8'd138;
		data_a[14374]<=8'd124;
		data_a[14375]<=8'd96;
		data_a[14376]<=8'd90;
		data_a[14377]<=8'd89;
		data_a[14378]<=8'd73;
		data_a[14379]<=8'd88;
		data_a[14380]<=8'd75;
		data_a[14381]<=8'd91;
		data_a[14382]<=8'd129;
		data_a[14383]<=8'd218;
		data_a[14384]<=8'd238;
		data_a[14385]<=8'd238;
		data_a[14386]<=8'd239;
		data_a[14387]<=8'd239;
		data_a[14388]<=8'd239;
		data_a[14389]<=8'd240;
		data_a[14390]<=8'd241;
		data_a[14391]<=8'd241;
		data_a[14392]<=8'd241;
		data_a[14393]<=8'd242;
		data_a[14394]<=8'd243;
		data_a[14395]<=8'd244;
		data_a[14396]<=8'd245;
		data_a[14397]<=8'd246;
		data_a[14398]<=8'd247;
		data_a[14399]<=8'd247;
		data_a[14400]<=8'd255;
		data_a[14401]<=8'd81;
		data_a[14402]<=8'd80;
		data_a[14403]<=8'd80;
		data_a[14404]<=8'd79;
		data_a[14405]<=8'd79;
		data_a[14406]<=8'd78;
		data_a[14407]<=8'd69;
		data_a[14408]<=8'd64;
		data_a[14409]<=8'd59;
		data_a[14410]<=8'd63;
		data_a[14411]<=8'd65;
		data_a[14412]<=8'd65;
		data_a[14413]<=8'd69;
		data_a[14414]<=8'd70;
		data_a[14415]<=8'd70;
		data_a[14416]<=8'd67;
		data_a[14417]<=8'd65;
		data_a[14418]<=8'd56;
		data_a[14419]<=8'd50;
		data_a[14420]<=8'd47;
		data_a[14421]<=8'd65;
		data_a[14422]<=8'd63;
		data_a[14423]<=8'd50;
		data_a[14424]<=8'd111;
		data_a[14425]<=8'd123;
		data_a[14426]<=8'd94;
		data_a[14427]<=8'd83;
		data_a[14428]<=8'd145;
		data_a[14429]<=8'd143;
		data_a[14430]<=8'd148;
		data_a[14431]<=8'd163;
		data_a[14432]<=8'd157;
		data_a[14433]<=8'd158;
		data_a[14434]<=8'd154;
		data_a[14435]<=8'd159;
		data_a[14436]<=8'd154;
		data_a[14437]<=8'd121;
		data_a[14438]<=8'd107;
		data_a[14439]<=8'd92;
		data_a[14440]<=8'd86;
		data_a[14441]<=8'd66;
		data_a[14442]<=8'd123;
		data_a[14443]<=8'd151;
		data_a[14444]<=8'd170;
		data_a[14445]<=8'd170;
		data_a[14446]<=8'd177;
		data_a[14447]<=8'd197;
		data_a[14448]<=8'd185;
		data_a[14449]<=8'd164;
		data_a[14450]<=8'd129;
		data_a[14451]<=8'd106;
		data_a[14452]<=8'd53;
		data_a[14453]<=8'd85;
		data_a[14454]<=8'd102;
		data_a[14455]<=8'd107;
		data_a[14456]<=8'd115;
		data_a[14457]<=8'd117;
		data_a[14458]<=8'd127;
		data_a[14459]<=8'd123;
		data_a[14460]<=8'd117;
		data_a[14461]<=8'd142;
		data_a[14462]<=8'd92;
		data_a[14463]<=8'd134;
		data_a[14464]<=8'd149;
		data_a[14465]<=8'd112;
		data_a[14466]<=8'd85;
		data_a[14467]<=8'd101;
		data_a[14468]<=8'd97;
		data_a[14469]<=8'd157;
		data_a[14470]<=8'd182;
		data_a[14471]<=8'd210;
		data_a[14472]<=8'd215;
		data_a[14473]<=8'd213;
		data_a[14474]<=8'd217;
		data_a[14475]<=8'd218;
		data_a[14476]<=8'd215;
		data_a[14477]<=8'd227;
		data_a[14478]<=8'd230;
		data_a[14479]<=8'd227;
		data_a[14480]<=8'd225;
		data_a[14481]<=8'd229;
		data_a[14482]<=8'd237;
		data_a[14483]<=8'd112;
		data_a[14484]<=8'd80;
		data_a[14485]<=8'd134;
		data_a[14486]<=8'd139;
		data_a[14487]<=8'd144;
		data_a[14488]<=8'd154;
		data_a[14489]<=8'd161;
		data_a[14490]<=8'd169;
		data_a[14491]<=8'd164;
		data_a[14492]<=8'd162;
		data_a[14493]<=8'd168;
		data_a[14494]<=8'd165;
		data_a[14495]<=8'd163;
		data_a[14496]<=8'd154;
		data_a[14497]<=8'd142;
		data_a[14498]<=8'd115;
		data_a[14499]<=8'd90;
		data_a[14500]<=8'd77;
		data_a[14501]<=8'd75;
		data_a[14502]<=8'd70;
		data_a[14503]<=8'd68;
		data_a[14504]<=8'd69;
		data_a[14505]<=8'd77;
		data_a[14506]<=8'd80;
		data_a[14507]<=8'd75;
		data_a[14508]<=8'd77;
		data_a[14509]<=8'd79;
		data_a[14510]<=8'd73;
		data_a[14511]<=8'd66;
		data_a[14512]<=8'd71;
		data_a[14513]<=8'd75;
		data_a[14514]<=8'd71;
		data_a[14515]<=8'd72;
		data_a[14516]<=8'd61;
		data_a[14517]<=8'd64;
		data_a[14518]<=8'd74;
		data_a[14519]<=8'd75;
		data_a[14520]<=8'd68;
		data_a[14521]<=8'd85;
		data_a[14522]<=8'd136;
		data_a[14523]<=8'd134;
		data_a[14524]<=8'd111;
		data_a[14525]<=8'd87;
		data_a[14526]<=8'd88;
		data_a[14527]<=8'd82;
		data_a[14528]<=8'd79;
		data_a[14529]<=8'd86;
		data_a[14530]<=8'd71;
		data_a[14531]<=8'd84;
		data_a[14532]<=8'd143;
		data_a[14533]<=8'd176;
		data_a[14534]<=8'd241;
		data_a[14535]<=8'd238;
		data_a[14536]<=8'd238;
		data_a[14537]<=8'd238;
		data_a[14538]<=8'd239;
		data_a[14539]<=8'd240;
		data_a[14540]<=8'd241;
		data_a[14541]<=8'd242;
		data_a[14542]<=8'd242;
		data_a[14543]<=8'd242;
		data_a[14544]<=8'd244;
		data_a[14545]<=8'd245;
		data_a[14546]<=8'd246;
		data_a[14547]<=8'd246;
		data_a[14548]<=8'd247;
		data_a[14549]<=8'd247;
		data_a[14550]<=8'd255;
		data_a[14551]<=8'd80;
		data_a[14552]<=8'd78;
		data_a[14553]<=8'd79;
		data_a[14554]<=8'd78;
		data_a[14555]<=8'd78;
		data_a[14556]<=8'd77;
		data_a[14557]<=8'd68;
		data_a[14558]<=8'd62;
		data_a[14559]<=8'd56;
		data_a[14560]<=8'd62;
		data_a[14561]<=8'd67;
		data_a[14562]<=8'd68;
		data_a[14563]<=8'd71;
		data_a[14564]<=8'd71;
		data_a[14565]<=8'd71;
		data_a[14566]<=8'd71;
		data_a[14567]<=8'd66;
		data_a[14568]<=8'd54;
		data_a[14569]<=8'd50;
		data_a[14570]<=8'd45;
		data_a[14571]<=8'd101;
		data_a[14572]<=8'd67;
		data_a[14573]<=8'd49;
		data_a[14574]<=8'd122;
		data_a[14575]<=8'd160;
		data_a[14576]<=8'd116;
		data_a[14577]<=8'd86;
		data_a[14578]<=8'd141;
		data_a[14579]<=8'd149;
		data_a[14580]<=8'd150;
		data_a[14581]<=8'd154;
		data_a[14582]<=8'd165;
		data_a[14583]<=8'd159;
		data_a[14584]<=8'd142;
		data_a[14585]<=8'd120;
		data_a[14586]<=8'd117;
		data_a[14587]<=8'd106;
		data_a[14588]<=8'd110;
		data_a[14589]<=8'd101;
		data_a[14590]<=8'd100;
		data_a[14591]<=8'd125;
		data_a[14592]<=8'd149;
		data_a[14593]<=8'd156;
		data_a[14594]<=8'd173;
		data_a[14595]<=8'd169;
		data_a[14596]<=8'd181;
		data_a[14597]<=8'd189;
		data_a[14598]<=8'd177;
		data_a[14599]<=8'd164;
		data_a[14600]<=8'd142;
		data_a[14601]<=8'd132;
		data_a[14602]<=8'd75;
		data_a[14603]<=8'd92;
		data_a[14604]<=8'd55;
		data_a[14605]<=8'd65;
		data_a[14606]<=8'd87;
		data_a[14607]<=8'd103;
		data_a[14608]<=8'd104;
		data_a[14609]<=8'd107;
		data_a[14610]<=8'd55;
		data_a[14611]<=8'd62;
		data_a[14612]<=8'd126;
		data_a[14613]<=8'd145;
		data_a[14614]<=8'd148;
		data_a[14615]<=8'd105;
		data_a[14616]<=8'd93;
		data_a[14617]<=8'd122;
		data_a[14618]<=8'd123;
		data_a[14619]<=8'd184;
		data_a[14620]<=8'd199;
		data_a[14621]<=8'd214;
		data_a[14622]<=8'd217;
		data_a[14623]<=8'd217;
		data_a[14624]<=8'd219;
		data_a[14625]<=8'd220;
		data_a[14626]<=8'd218;
		data_a[14627]<=8'd229;
		data_a[14628]<=8'd229;
		data_a[14629]<=8'd228;
		data_a[14630]<=8'd231;
		data_a[14631]<=8'd228;
		data_a[14632]<=8'd221;
		data_a[14633]<=8'd128;
		data_a[14634]<=8'd70;
		data_a[14635]<=8'd130;
		data_a[14636]<=8'd141;
		data_a[14637]<=8'd138;
		data_a[14638]<=8'd158;
		data_a[14639]<=8'd162;
		data_a[14640]<=8'd167;
		data_a[14641]<=8'd156;
		data_a[14642]<=8'd161;
		data_a[14643]<=8'd156;
		data_a[14644]<=8'd160;
		data_a[14645]<=8'd145;
		data_a[14646]<=8'd130;
		data_a[14647]<=8'd122;
		data_a[14648]<=8'd89;
		data_a[14649]<=8'd76;
		data_a[14650]<=8'd80;
		data_a[14651]<=8'd78;
		data_a[14652]<=8'd66;
		data_a[14653]<=8'd75;
		data_a[14654]<=8'd69;
		data_a[14655]<=8'd99;
		data_a[14656]<=8'd109;
		data_a[14657]<=8'd88;
		data_a[14658]<=8'd78;
		data_a[14659]<=8'd84;
		data_a[14660]<=8'd67;
		data_a[14661]<=8'd68;
		data_a[14662]<=8'd60;
		data_a[14663]<=8'd67;
		data_a[14664]<=8'd71;
		data_a[14665]<=8'd65;
		data_a[14666]<=8'd57;
		data_a[14667]<=8'd61;
		data_a[14668]<=8'd73;
		data_a[14669]<=8'd74;
		data_a[14670]<=8'd67;
		data_a[14671]<=8'd85;
		data_a[14672]<=8'd137;
		data_a[14673]<=8'd129;
		data_a[14674]<=8'd105;
		data_a[14675]<=8'd83;
		data_a[14676]<=8'd81;
		data_a[14677]<=8'd81;
		data_a[14678]<=8'd86;
		data_a[14679]<=8'd72;
		data_a[14680]<=8'd75;
		data_a[14681]<=8'd83;
		data_a[14682]<=8'd181;
		data_a[14683]<=8'd185;
		data_a[14684]<=8'd234;
		data_a[14685]<=8'd235;
		data_a[14686]<=8'd239;
		data_a[14687]<=8'd240;
		data_a[14688]<=8'd240;
		data_a[14689]<=8'd240;
		data_a[14690]<=8'd240;
		data_a[14691]<=8'd241;
		data_a[14692]<=8'd242;
		data_a[14693]<=8'd243;
		data_a[14694]<=8'd244;
		data_a[14695]<=8'd245;
		data_a[14696]<=8'd246;
		data_a[14697]<=8'd246;
		data_a[14698]<=8'd247;
		data_a[14699]<=8'd247;
		data_a[14700]<=8'd255;
		data_a[14701]<=8'd77;
		data_a[14702]<=8'd75;
		data_a[14703]<=8'd77;
		data_a[14704]<=8'd77;
		data_a[14705]<=8'd76;
		data_a[14706]<=8'd75;
		data_a[14707]<=8'd67;
		data_a[14708]<=8'd63;
		data_a[14709]<=8'd57;
		data_a[14710]<=8'd64;
		data_a[14711]<=8'd72;
		data_a[14712]<=8'd73;
		data_a[14713]<=8'd72;
		data_a[14714]<=8'd70;
		data_a[14715]<=8'd69;
		data_a[14716]<=8'd63;
		data_a[14717]<=8'd66;
		data_a[14718]<=8'd57;
		data_a[14719]<=8'd53;
		data_a[14720]<=8'd45;
		data_a[14721]<=8'd142;
		data_a[14722]<=8'd119;
		data_a[14723]<=8'd120;
		data_a[14724]<=8'd143;
		data_a[14725]<=8'd150;
		data_a[14726]<=8'd128;
		data_a[14727]<=8'd95;
		data_a[14728]<=8'd134;
		data_a[14729]<=8'd146;
		data_a[14730]<=8'd151;
		data_a[14731]<=8'd156;
		data_a[14732]<=8'd161;
		data_a[14733]<=8'd157;
		data_a[14734]<=8'd152;
		data_a[14735]<=8'd133;
		data_a[14736]<=8'd136;
		data_a[14737]<=8'd126;
		data_a[14738]<=8'd127;
		data_a[14739]<=8'd119;
		data_a[14740]<=8'd136;
		data_a[14741]<=8'd124;
		data_a[14742]<=8'd134;
		data_a[14743]<=8'd149;
		data_a[14744]<=8'd166;
		data_a[14745]<=8'd169;
		data_a[14746]<=8'd177;
		data_a[14747]<=8'd186;
		data_a[14748]<=8'd181;
		data_a[14749]<=8'd154;
		data_a[14750]<=8'd135;
		data_a[14751]<=8'd132;
		data_a[14752]<=8'd121;
		data_a[14753]<=8'd97;
		data_a[14754]<=8'd115;
		data_a[14755]<=8'd114;
		data_a[14756]<=8'd114;
		data_a[14757]<=8'd119;
		data_a[14758]<=8'd116;
		data_a[14759]<=8'd114;
		data_a[14760]<=8'd125;
		data_a[14761]<=8'd138;
		data_a[14762]<=8'd141;
		data_a[14763]<=8'd147;
		data_a[14764]<=8'd133;
		data_a[14765]<=8'd97;
		data_a[14766]<=8'd110;
		data_a[14767]<=8'd110;
		data_a[14768]<=8'd119;
		data_a[14769]<=8'd128;
		data_a[14770]<=8'd215;
		data_a[14771]<=8'd224;
		data_a[14772]<=8'd218;
		data_a[14773]<=8'd221;
		data_a[14774]<=8'd221;
		data_a[14775]<=8'd221;
		data_a[14776]<=8'd220;
		data_a[14777]<=8'd230;
		data_a[14778]<=8'd229;
		data_a[14779]<=8'd229;
		data_a[14780]<=8'd228;
		data_a[14781]<=8'd227;
		data_a[14782]<=8'd222;
		data_a[14783]<=8'd223;
		data_a[14784]<=8'd79;
		data_a[14785]<=8'd120;
		data_a[14786]<=8'd127;
		data_a[14787]<=8'd145;
		data_a[14788]<=8'd149;
		data_a[14789]<=8'd160;
		data_a[14790]<=8'd155;
		data_a[14791]<=8'd159;
		data_a[14792]<=8'd152;
		data_a[14793]<=8'd148;
		data_a[14794]<=8'd138;
		data_a[14795]<=8'd111;
		data_a[14796]<=8'd102;
		data_a[14797]<=8'd97;
		data_a[14798]<=8'd79;
		data_a[14799]<=8'd77;
		data_a[14800]<=8'd69;
		data_a[14801]<=8'd71;
		data_a[14802]<=8'd66;
		data_a[14803]<=8'd72;
		data_a[14804]<=8'd85;
		data_a[14805]<=8'd105;
		data_a[14806]<=8'd108;
		data_a[14807]<=8'd97;
		data_a[14808]<=8'd78;
		data_a[14809]<=8'd85;
		data_a[14810]<=8'd78;
		data_a[14811]<=8'd72;
		data_a[14812]<=8'd60;
		data_a[14813]<=8'd66;
		data_a[14814]<=8'd75;
		data_a[14815]<=8'd63;
		data_a[14816]<=8'd61;
		data_a[14817]<=8'd69;
		data_a[14818]<=8'd79;
		data_a[14819]<=8'd76;
		data_a[14820]<=8'd74;
		data_a[14821]<=8'd90;
		data_a[14822]<=8'd136;
		data_a[14823]<=8'd123;
		data_a[14824]<=8'd100;
		data_a[14825]<=8'd82;
		data_a[14826]<=8'd75;
		data_a[14827]<=8'd78;
		data_a[14828]<=8'd81;
		data_a[14829]<=8'd81;
		data_a[14830]<=8'd78;
		data_a[14831]<=8'd79;
		data_a[14832]<=8'd120;
		data_a[14833]<=8'd222;
		data_a[14834]<=8'd239;
		data_a[14835]<=8'd245;
		data_a[14836]<=8'd240;
		data_a[14837]<=8'd241;
		data_a[14838]<=8'd241;
		data_a[14839]<=8'd241;
		data_a[14840]<=8'd240;
		data_a[14841]<=8'd241;
		data_a[14842]<=8'd242;
		data_a[14843]<=8'd244;
		data_a[14844]<=8'd245;
		data_a[14845]<=8'd245;
		data_a[14846]<=8'd246;
		data_a[14847]<=8'd246;
		data_a[14848]<=8'd247;
		data_a[14849]<=8'd247;
		data_a[14850]<=8'd254;
		data_a[14851]<=8'd76;
		data_a[14852]<=8'd74;
		data_a[14853]<=8'd77;
		data_a[14854]<=8'd77;
		data_a[14855]<=8'd75;
		data_a[14856]<=8'd74;
		data_a[14857]<=8'd67;
		data_a[14858]<=8'd65;
		data_a[14859]<=8'd57;
		data_a[14860]<=8'd65;
		data_a[14861]<=8'd74;
		data_a[14862]<=8'd75;
		data_a[14863]<=8'd72;
		data_a[14864]<=8'd68;
		data_a[14865]<=8'd69;
		data_a[14866]<=8'd68;
		data_a[14867]<=8'd67;
		data_a[14868]<=8'd53;
		data_a[14869]<=8'd50;
		data_a[14870]<=8'd44;
		data_a[14871]<=8'd145;
		data_a[14872]<=8'd128;
		data_a[14873]<=8'd129;
		data_a[14874]<=8'd176;
		data_a[14875]<=8'd129;
		data_a[14876]<=8'd140;
		data_a[14877]<=8'd92;
		data_a[14878]<=8'd125;
		data_a[14879]<=8'd147;
		data_a[14880]<=8'd142;
		data_a[14881]<=8'd157;
		data_a[14882]<=8'd150;
		data_a[14883]<=8'd144;
		data_a[14884]<=8'd144;
		data_a[14885]<=8'd133;
		data_a[14886]<=8'd138;
		data_a[14887]<=8'd134;
		data_a[14888]<=8'd129;
		data_a[14889]<=8'd126;
		data_a[14890]<=8'd116;
		data_a[14891]<=8'd109;
		data_a[14892]<=8'd145;
		data_a[14893]<=8'd165;
		data_a[14894]<=8'd160;
		data_a[14895]<=8'd156;
		data_a[14896]<=8'd178;
		data_a[14897]<=8'd183;
		data_a[14898]<=8'd162;
		data_a[14899]<=8'd154;
		data_a[14900]<=8'd142;
		data_a[14901]<=8'd130;
		data_a[14902]<=8'd117;
		data_a[14903]<=8'd119;
		data_a[14904]<=8'd101;
		data_a[14905]<=8'd113;
		data_a[14906]<=8'd109;
		data_a[14907]<=8'd115;
		data_a[14908]<=8'd107;
		data_a[14909]<=8'd115;
		data_a[14910]<=8'd124;
		data_a[14911]<=8'd137;
		data_a[14912]<=8'd146;
		data_a[14913]<=8'd144;
		data_a[14914]<=8'd117;
		data_a[14915]<=8'd116;
		data_a[14916]<=8'd129;
		data_a[14917]<=8'd79;
		data_a[14918]<=8'd102;
		data_a[14919]<=8'd215;
		data_a[14920]<=8'd213;
		data_a[14921]<=8'd218;
		data_a[14922]<=8'd218;
		data_a[14923]<=8'd222;
		data_a[14924]<=8'd222;
		data_a[14925]<=8'd220;
		data_a[14926]<=8'd221;
		data_a[14927]<=8'd231;
		data_a[14928]<=8'd229;
		data_a[14929]<=8'd230;
		data_a[14930]<=8'd232;
		data_a[14931]<=8'd234;
		data_a[14932]<=8'd223;
		data_a[14933]<=8'd203;
		data_a[14934]<=8'd83;
		data_a[14935]<=8'd97;
		data_a[14936]<=8'd130;
		data_a[14937]<=8'd131;
		data_a[14938]<=8'd151;
		data_a[14939]<=8'd155;
		data_a[14940]<=8'd154;
		data_a[14941]<=8'd149;
		data_a[14942]<=8'd148;
		data_a[14943]<=8'd134;
		data_a[14944]<=8'd124;
		data_a[14945]<=8'd91;
		data_a[14946]<=8'd90;
		data_a[14947]<=8'd77;
		data_a[14948]<=8'd72;
		data_a[14949]<=8'd87;
		data_a[14950]<=8'd70;
		data_a[14951]<=8'd68;
		data_a[14952]<=8'd61;
		data_a[14953]<=8'd61;
		data_a[14954]<=8'd89;
		data_a[14955]<=8'd89;
		data_a[14956]<=8'd108;
		data_a[14957]<=8'd100;
		data_a[14958]<=8'd80;
		data_a[14959]<=8'd86;
		data_a[14960]<=8'd67;
		data_a[14961]<=8'd64;
		data_a[14962]<=8'd76;
		data_a[14963]<=8'd77;
		data_a[14964]<=8'd86;
		data_a[14965]<=8'd80;
		data_a[14966]<=8'd81;
		data_a[14967]<=8'd88;
		data_a[14968]<=8'd84;
		data_a[14969]<=8'd72;
		data_a[14970]<=8'd79;
		data_a[14971]<=8'd96;
		data_a[14972]<=8'd128;
		data_a[14973]<=8'd114;
		data_a[14974]<=8'd97;
		data_a[14975]<=8'd80;
		data_a[14976]<=8'd74;
		data_a[14977]<=8'd74;
		data_a[14978]<=8'd71;
		data_a[14979]<=8'd71;
		data_a[14980]<=8'd73;
		data_a[14981]<=8'd91;
		data_a[14982]<=8'd111;
		data_a[14983]<=8'd226;
		data_a[14984]<=8'd245;
		data_a[14985]<=8'd243;
		data_a[14986]<=8'd240;
		data_a[14987]<=8'd241;
		data_a[14988]<=8'd242;
		data_a[14989]<=8'd242;
		data_a[14990]<=8'd242;
		data_a[14991]<=8'd242;
		data_a[14992]<=8'd244;
		data_a[14993]<=8'd245;
		data_a[14994]<=8'd245;
		data_a[14995]<=8'd245;
		data_a[14996]<=8'd246;
		data_a[14997]<=8'd247;
		data_a[14998]<=8'd247;
		data_a[14999]<=8'd248;
		data_a[15000]<=8'd255;
		data_a[15001]<=8'd78;
		data_a[15002]<=8'd77;
		data_a[15003]<=8'd80;
		data_a[15004]<=8'd79;
		data_a[15005]<=8'd77;
		data_a[15006]<=8'd76;
		data_a[15007]<=8'd68;
		data_a[15008]<=8'd64;
		data_a[15009]<=8'd56;
		data_a[15010]<=8'd63;
		data_a[15011]<=8'd73;
		data_a[15012]<=8'd73;
		data_a[15013]<=8'd70;
		data_a[15014]<=8'd67;
		data_a[15015]<=8'd69;
		data_a[15016]<=8'd70;
		data_a[15017]<=8'd65;
		data_a[15018]<=8'd54;
		data_a[15019]<=8'd54;
		data_a[15020]<=8'd52;
		data_a[15021]<=8'd156;
		data_a[15022]<=8'd132;
		data_a[15023]<=8'd129;
		data_a[15024]<=8'd154;
		data_a[15025]<=8'd166;
		data_a[15026]<=8'd154;
		data_a[15027]<=8'd95;
		data_a[15028]<=8'd127;
		data_a[15029]<=8'd142;
		data_a[15030]<=8'd156;
		data_a[15031]<=8'd143;
		data_a[15032]<=8'd139;
		data_a[15033]<=8'd140;
		data_a[15034]<=8'd143;
		data_a[15035]<=8'd136;
		data_a[15036]<=8'd135;
		data_a[15037]<=8'd133;
		data_a[15038]<=8'd115;
		data_a[15039]<=8'd106;
		data_a[15040]<=8'd102;
		data_a[15041]<=8'd108;
		data_a[15042]<=8'd169;
		data_a[15043]<=8'd167;
		data_a[15044]<=8'd172;
		data_a[15045]<=8'd175;
		data_a[15046]<=8'd165;
		data_a[15047]<=8'd166;
		data_a[15048]<=8'd154;
		data_a[15049]<=8'd150;
		data_a[15050]<=8'd148;
		data_a[15051]<=8'd143;
		data_a[15052]<=8'd119;
		data_a[15053]<=8'd99;
		data_a[15054]<=8'd112;
		data_a[15055]<=8'd109;
		data_a[15056]<=8'd107;
		data_a[15057]<=8'd110;
		data_a[15058]<=8'd108;
		data_a[15059]<=8'd107;
		data_a[15060]<=8'd126;
		data_a[15061]<=8'd140;
		data_a[15062]<=8'd137;
		data_a[15063]<=8'd150;
		data_a[15064]<=8'd93;
		data_a[15065]<=8'd128;
		data_a[15066]<=8'd129;
		data_a[15067]<=8'd81;
		data_a[15068]<=8'd108;
		data_a[15069]<=8'd194;
		data_a[15070]<=8'd220;
		data_a[15071]<=8'd221;
		data_a[15072]<=8'd219;
		data_a[15073]<=8'd223;
		data_a[15074]<=8'd222;
		data_a[15075]<=8'd219;
		data_a[15076]<=8'd221;
		data_a[15077]<=8'd232;
		data_a[15078]<=8'd231;
		data_a[15079]<=8'd232;
		data_a[15080]<=8'd231;
		data_a[15081]<=8'd232;
		data_a[15082]<=8'd226;
		data_a[15083]<=8'd215;
		data_a[15084]<=8'd84;
		data_a[15085]<=8'd77;
		data_a[15086]<=8'd121;
		data_a[15087]<=8'd131;
		data_a[15088]<=8'd149;
		data_a[15089]<=8'd151;
		data_a[15090]<=8'd153;
		data_a[15091]<=8'd145;
		data_a[15092]<=8'd142;
		data_a[15093]<=8'd125;
		data_a[15094]<=8'd107;
		data_a[15095]<=8'd78;
		data_a[15096]<=8'd79;
		data_a[15097]<=8'd67;
		data_a[15098]<=8'd68;
		data_a[15099]<=8'd91;
		data_a[15100]<=8'd75;
		data_a[15101]<=8'd65;
		data_a[15102]<=8'd57;
		data_a[15103]<=8'd68;
		data_a[15104]<=8'd87;
		data_a[15105]<=8'd94;
		data_a[15106]<=8'd95;
		data_a[15107]<=8'd92;
		data_a[15108]<=8'd84;
		data_a[15109]<=8'd76;
		data_a[15110]<=8'd79;
		data_a[15111]<=8'd90;
		data_a[15112]<=8'd101;
		data_a[15113]<=8'd95;
		data_a[15114]<=8'd94;
		data_a[15115]<=8'd93;
		data_a[15116]<=8'd93;
		data_a[15117]<=8'd101;
		data_a[15118]<=8'd90;
		data_a[15119]<=8'd77;
		data_a[15120]<=8'd76;
		data_a[15121]<=8'd97;
		data_a[15122]<=8'd117;
		data_a[15123]<=8'd109;
		data_a[15124]<=8'd92;
		data_a[15125]<=8'd72;
		data_a[15126]<=8'd73;
		data_a[15127]<=8'd69;
		data_a[15128]<=8'd70;
		data_a[15129]<=8'd74;
		data_a[15130]<=8'd72;
		data_a[15131]<=8'd81;
		data_a[15132]<=8'd119;
		data_a[15133]<=8'd253;
		data_a[15134]<=8'd241;
		data_a[15135]<=8'd240;
		data_a[15136]<=8'd241;
		data_a[15137]<=8'd241;
		data_a[15138]<=8'd242;
		data_a[15139]<=8'd243;
		data_a[15140]<=8'd244;
		data_a[15141]<=8'd244;
		data_a[15142]<=8'd244;
		data_a[15143]<=8'd244;
		data_a[15144]<=8'd245;
		data_a[15145]<=8'd246;
		data_a[15146]<=8'd246;
		data_a[15147]<=8'd247;
		data_a[15148]<=8'd247;
		data_a[15149]<=8'd248;
		data_a[15150]<=8'd254;
		data_a[15151]<=8'd79;
		data_a[15152]<=8'd80;
		data_a[15153]<=8'd81;
		data_a[15154]<=8'd80;
		data_a[15155]<=8'd78;
		data_a[15156]<=8'd76;
		data_a[15157]<=8'd67;
		data_a[15158]<=8'd66;
		data_a[15159]<=8'd59;
		data_a[15160]<=8'd65;
		data_a[15161]<=8'd73;
		data_a[15162]<=8'd71;
		data_a[15163]<=8'd69;
		data_a[15164]<=8'd68;
		data_a[15165]<=8'd70;
		data_a[15166]<=8'd67;
		data_a[15167]<=8'd64;
		data_a[15168]<=8'd59;
		data_a[15169]<=8'd57;
		data_a[15170]<=8'd46;
		data_a[15171]<=8'd161;
		data_a[15172]<=8'd131;
		data_a[15173]<=8'd133;
		data_a[15174]<=8'd138;
		data_a[15175]<=8'd155;
		data_a[15176]<=8'd138;
		data_a[15177]<=8'd88;
		data_a[15178]<=8'd122;
		data_a[15179]<=8'd143;
		data_a[15180]<=8'd143;
		data_a[15181]<=8'd144;
		data_a[15182]<=8'd140;
		data_a[15183]<=8'd137;
		data_a[15184]<=8'd134;
		data_a[15185]<=8'd132;
		data_a[15186]<=8'd125;
		data_a[15187]<=8'd117;
		data_a[15188]<=8'd100;
		data_a[15189]<=8'd99;
		data_a[15190]<=8'd101;
		data_a[15191]<=8'd121;
		data_a[15192]<=8'd162;
		data_a[15193]<=8'd165;
		data_a[15194]<=8'd175;
		data_a[15195]<=8'd166;
		data_a[15196]<=8'd166;
		data_a[15197]<=8'd152;
		data_a[15198]<=8'd144;
		data_a[15199]<=8'd142;
		data_a[15200]<=8'd153;
		data_a[15201]<=8'd153;
		data_a[15202]<=8'd144;
		data_a[15203]<=8'd87;
		data_a[15204]<=8'd102;
		data_a[15205]<=8'd125;
		data_a[15206]<=8'd122;
		data_a[15207]<=8'd118;
		data_a[15208]<=8'd117;
		data_a[15209]<=8'd114;
		data_a[15210]<=8'd133;
		data_a[15211]<=8'd142;
		data_a[15212]<=8'd143;
		data_a[15213]<=8'd152;
		data_a[15214]<=8'd85;
		data_a[15215]<=8'd108;
		data_a[15216]<=8'd121;
		data_a[15217]<=8'd65;
		data_a[15218]<=8'd123;
		data_a[15219]<=8'd225;
		data_a[15220]<=8'd229;
		data_a[15221]<=8'd223;
		data_a[15222]<=8'd221;
		data_a[15223]<=8'd224;
		data_a[15224]<=8'd223;
		data_a[15225]<=8'd221;
		data_a[15226]<=8'd221;
		data_a[15227]<=8'd233;
		data_a[15228]<=8'd234;
		data_a[15229]<=8'd234;
		data_a[15230]<=8'd230;
		data_a[15231]<=8'd238;
		data_a[15232]<=8'd223;
		data_a[15233]<=8'd190;
		data_a[15234]<=8'd87;
		data_a[15235]<=8'd75;
		data_a[15236]<=8'd109;
		data_a[15237]<=8'd126;
		data_a[15238]<=8'd141;
		data_a[15239]<=8'd149;
		data_a[15240]<=8'd148;
		data_a[15241]<=8'd148;
		data_a[15242]<=8'd133;
		data_a[15243]<=8'd114;
		data_a[15244]<=8'd87;
		data_a[15245]<=8'd69;
		data_a[15246]<=8'd67;
		data_a[15247]<=8'd66;
		data_a[15248]<=8'd74;
		data_a[15249]<=8'd88;
		data_a[15250]<=8'd68;
		data_a[15251]<=8'd67;
		data_a[15252]<=8'd69;
		data_a[15253]<=8'd75;
		data_a[15254]<=8'd88;
		data_a[15255]<=8'd94;
		data_a[15256]<=8'd97;
		data_a[15257]<=8'd76;
		data_a[15258]<=8'd79;
		data_a[15259]<=8'd102;
		data_a[15260]<=8'd107;
		data_a[15261]<=8'd108;
		data_a[15262]<=8'd110;
		data_a[15263]<=8'd104;
		data_a[15264]<=8'd101;
		data_a[15265]<=8'd105;
		data_a[15266]<=8'd105;
		data_a[15267]<=8'd112;
		data_a[15268]<=8'd103;
		data_a[15269]<=8'd93;
		data_a[15270]<=8'd77;
		data_a[15271]<=8'd101;
		data_a[15272]<=8'd115;
		data_a[15273]<=8'd110;
		data_a[15274]<=8'd89;
		data_a[15275]<=8'd64;
		data_a[15276]<=8'd70;
		data_a[15277]<=8'd66;
		data_a[15278]<=8'd64;
		data_a[15279]<=8'd76;
		data_a[15280]<=8'd68;
		data_a[15281]<=8'd78;
		data_a[15282]<=8'd138;
		data_a[15283]<=8'd239;
		data_a[15284]<=8'd243;
		data_a[15285]<=8'd236;
		data_a[15286]<=8'd243;
		data_a[15287]<=8'd243;
		data_a[15288]<=8'd243;
		data_a[15289]<=8'd244;
		data_a[15290]<=8'd245;
		data_a[15291]<=8'd245;
		data_a[15292]<=8'd244;
		data_a[15293]<=8'd243;
		data_a[15294]<=8'd246;
		data_a[15295]<=8'd246;
		data_a[15296]<=8'd246;
		data_a[15297]<=8'd247;
		data_a[15298]<=8'd247;
		data_a[15299]<=8'd248;
		data_a[15300]<=8'd254;
		data_a[15301]<=8'd81;
		data_a[15302]<=8'd81;
		data_a[15303]<=8'd82;
		data_a[15304]<=8'd80;
		data_a[15305]<=8'd80;
		data_a[15306]<=8'd76;
		data_a[15307]<=8'd63;
		data_a[15308]<=8'd69;
		data_a[15309]<=8'd62;
		data_a[15310]<=8'd69;
		data_a[15311]<=8'd74;
		data_a[15312]<=8'd71;
		data_a[15313]<=8'd69;
		data_a[15314]<=8'd69;
		data_a[15315]<=8'd71;
		data_a[15316]<=8'd66;
		data_a[15317]<=8'd63;
		data_a[15318]<=8'd56;
		data_a[15319]<=8'd60;
		data_a[15320]<=8'd50;
		data_a[15321]<=8'd161;
		data_a[15322]<=8'd134;
		data_a[15323]<=8'd132;
		data_a[15324]<=8'd99;
		data_a[15325]<=8'd125;
		data_a[15326]<=8'd127;
		data_a[15327]<=8'd93;
		data_a[15328]<=8'd120;
		data_a[15329]<=8'd145;
		data_a[15330]<=8'd144;
		data_a[15331]<=8'd134;
		data_a[15332]<=8'd137;
		data_a[15333]<=8'd131;
		data_a[15334]<=8'd128;
		data_a[15335]<=8'd129;
		data_a[15336]<=8'd120;
		data_a[15337]<=8'd104;
		data_a[15338]<=8'd96;
		data_a[15339]<=8'd104;
		data_a[15340]<=8'd107;
		data_a[15341]<=8'd112;
		data_a[15342]<=8'd149;
		data_a[15343]<=8'd149;
		data_a[15344]<=8'd154;
		data_a[15345]<=8'd160;
		data_a[15346]<=8'd158;
		data_a[15347]<=8'd136;
		data_a[15348]<=8'd133;
		data_a[15349]<=8'd129;
		data_a[15350]<=8'd149;
		data_a[15351]<=8'd143;
		data_a[15352]<=8'd141;
		data_a[15353]<=8'd83;
		data_a[15354]<=8'd98;
		data_a[15355]<=8'd114;
		data_a[15356]<=8'd122;
		data_a[15357]<=8'd125;
		data_a[15358]<=8'd124;
		data_a[15359]<=8'd124;
		data_a[15360]<=8'd130;
		data_a[15361]<=8'd138;
		data_a[15362]<=8'd142;
		data_a[15363]<=8'd156;
		data_a[15364]<=8'd99;
		data_a[15365]<=8'd100;
		data_a[15366]<=8'd128;
		data_a[15367]<=8'd100;
		data_a[15368]<=8'd212;
		data_a[15369]<=8'd216;
		data_a[15370]<=8'd217;
		data_a[15371]<=8'd224;
		data_a[15372]<=8'd224;
		data_a[15373]<=8'd225;
		data_a[15374]<=8'd226;
		data_a[15375]<=8'd224;
		data_a[15376]<=8'd222;
		data_a[15377]<=8'd234;
		data_a[15378]<=8'd236;
		data_a[15379]<=8'd233;
		data_a[15380]<=8'd238;
		data_a[15381]<=8'd233;
		data_a[15382]<=8'd230;
		data_a[15383]<=8'd190;
		data_a[15384]<=8'd79;
		data_a[15385]<=8'd71;
		data_a[15386]<=8'd102;
		data_a[15387]<=8'd120;
		data_a[15388]<=8'd142;
		data_a[15389]<=8'd148;
		data_a[15390]<=8'd147;
		data_a[15391]<=8'd137;
		data_a[15392]<=8'd130;
		data_a[15393]<=8'd92;
		data_a[15394]<=8'd83;
		data_a[15395]<=8'd72;
		data_a[15396]<=8'd67;
		data_a[15397]<=8'd67;
		data_a[15398]<=8'd72;
		data_a[15399]<=8'd77;
		data_a[15400]<=8'd68;
		data_a[15401]<=8'd74;
		data_a[15402]<=8'd74;
		data_a[15403]<=8'd67;
		data_a[15404]<=8'd74;
		data_a[15405]<=8'd77;
		data_a[15406]<=8'd82;
		data_a[15407]<=8'd108;
		data_a[15408]<=8'd118;
		data_a[15409]<=8'd119;
		data_a[15410]<=8'd124;
		data_a[15411]<=8'd120;
		data_a[15412]<=8'd110;
		data_a[15413]<=8'd111;
		data_a[15414]<=8'd116;
		data_a[15415]<=8'd125;
		data_a[15416]<=8'd126;
		data_a[15417]<=8'd123;
		data_a[15418]<=8'd111;
		data_a[15419]<=8'd93;
		data_a[15420]<=8'd85;
		data_a[15421]<=8'd103;
		data_a[15422]<=8'd116;
		data_a[15423]<=8'd109;
		data_a[15424]<=8'd84;
		data_a[15425]<=8'd62;
		data_a[15426]<=8'd68;
		data_a[15427]<=8'd67;
		data_a[15428]<=8'd63;
		data_a[15429]<=8'd68;
		data_a[15430]<=8'd74;
		data_a[15431]<=8'd78;
		data_a[15432]<=8'd121;
		data_a[15433]<=8'd229;
		data_a[15434]<=8'd241;
		data_a[15435]<=8'd242;
		data_a[15436]<=8'd244;
		data_a[15437]<=8'd244;
		data_a[15438]<=8'd244;
		data_a[15439]<=8'd244;
		data_a[15440]<=8'd244;
		data_a[15441]<=8'd244;
		data_a[15442]<=8'd245;
		data_a[15443]<=8'd245;
		data_a[15444]<=8'd246;
		data_a[15445]<=8'd246;
		data_a[15446]<=8'd247;
		data_a[15447]<=8'd247;
		data_a[15448]<=8'd247;
		data_a[15449]<=8'd247;
		data_a[15450]<=8'd255;
		data_a[15451]<=8'd83;
		data_a[15452]<=8'd83;
		data_a[15453]<=8'd83;
		data_a[15454]<=8'd82;
		data_a[15455]<=8'd81;
		data_a[15456]<=8'd76;
		data_a[15457]<=8'd61;
		data_a[15458]<=8'd66;
		data_a[15459]<=8'd62;
		data_a[15460]<=8'd69;
		data_a[15461]<=8'd73;
		data_a[15462]<=8'd71;
		data_a[15463]<=8'd70;
		data_a[15464]<=8'd71;
		data_a[15465]<=8'd73;
		data_a[15466]<=8'd67;
		data_a[15467]<=8'd68;
		data_a[15468]<=8'd53;
		data_a[15469]<=8'd61;
		data_a[15470]<=8'd51;
		data_a[15471]<=8'd148;
		data_a[15472]<=8'd142;
		data_a[15473]<=8'd141;
		data_a[15474]<=8'd99;
		data_a[15475]<=8'd66;
		data_a[15476]<=8'd55;
		data_a[15477]<=8'd52;
		data_a[15478]<=8'd116;
		data_a[15479]<=8'd139;
		data_a[15480]<=8'd134;
		data_a[15481]<=8'd131;
		data_a[15482]<=8'd133;
		data_a[15483]<=8'd131;
		data_a[15484]<=8'd126;
		data_a[15485]<=8'd116;
		data_a[15486]<=8'd106;
		data_a[15487]<=8'd96;
		data_a[15488]<=8'd99;
		data_a[15489]<=8'd107;
		data_a[15490]<=8'd116;
		data_a[15491]<=8'd106;
		data_a[15492]<=8'd129;
		data_a[15493]<=8'd134;
		data_a[15494]<=8'd131;
		data_a[15495]<=8'd132;
		data_a[15496]<=8'd136;
		data_a[15497]<=8'd131;
		data_a[15498]<=8'd124;
		data_a[15499]<=8'd127;
		data_a[15500]<=8'd121;
		data_a[15501]<=8'd127;
		data_a[15502]<=8'd132;
		data_a[15503]<=8'd81;
		data_a[15504]<=8'd87;
		data_a[15505]<=8'd110;
		data_a[15506]<=8'd114;
		data_a[15507]<=8'd126;
		data_a[15508]<=8'd112;
		data_a[15509]<=8'd126;
		data_a[15510]<=8'd128;
		data_a[15511]<=8'd144;
		data_a[15512]<=8'd146;
		data_a[15513]<=8'd156;
		data_a[15514]<=8'd102;
		data_a[15515]<=8'd119;
		data_a[15516]<=8'd124;
		data_a[15517]<=8'd174;
		data_a[15518]<=8'd214;
		data_a[15519]<=8'd221;
		data_a[15520]<=8'd229;
		data_a[15521]<=8'd224;
		data_a[15522]<=8'd226;
		data_a[15523]<=8'd225;
		data_a[15524]<=8'd228;
		data_a[15525]<=8'd226;
		data_a[15526]<=8'd222;
		data_a[15527]<=8'd235;
		data_a[15528]<=8'd236;
		data_a[15529]<=8'd231;
		data_a[15530]<=8'd235;
		data_a[15531]<=8'd233;
		data_a[15532]<=8'd243;
		data_a[15533]<=8'd211;
		data_a[15534]<=8'd89;
		data_a[15535]<=8'd71;
		data_a[15536]<=8'd86;
		data_a[15537]<=8'd115;
		data_a[15538]<=8'd130;
		data_a[15539]<=8'd146;
		data_a[15540]<=8'd137;
		data_a[15541]<=8'd139;
		data_a[15542]<=8'd123;
		data_a[15543]<=8'd83;
		data_a[15544]<=8'd73;
		data_a[15545]<=8'd68;
		data_a[15546]<=8'd61;
		data_a[15547]<=8'd70;
		data_a[15548]<=8'd69;
		data_a[15549]<=8'd73;
		data_a[15550]<=8'd76;
		data_a[15551]<=8'd66;
		data_a[15552]<=8'd56;
		data_a[15553]<=8'd70;
		data_a[15554]<=8'd90;
		data_a[15555]<=8'd120;
		data_a[15556]<=8'd119;
		data_a[15557]<=8'd121;
		data_a[15558]<=8'd122;
		data_a[15559]<=8'd127;
		data_a[15560]<=8'd120;
		data_a[15561]<=8'd117;
		data_a[15562]<=8'd127;
		data_a[15563]<=8'd126;
		data_a[15564]<=8'd127;
		data_a[15565]<=8'd130;
		data_a[15566]<=8'd133;
		data_a[15567]<=8'd124;
		data_a[15568]<=8'd114;
		data_a[15569]<=8'd90;
		data_a[15570]<=8'd90;
		data_a[15571]<=8'd98;
		data_a[15572]<=8'd110;
		data_a[15573]<=8'd101;
		data_a[15574]<=8'd78;
		data_a[15575]<=8'd62;
		data_a[15576]<=8'd67;
		data_a[15577]<=8'd68;
		data_a[15578]<=8'd65;
		data_a[15579]<=8'd68;
		data_a[15580]<=8'd68;
		data_a[15581]<=8'd84;
		data_a[15582]<=8'd120;
		data_a[15583]<=8'd230;
		data_a[15584]<=8'd242;
		data_a[15585]<=8'd243;
		data_a[15586]<=8'd244;
		data_a[15587]<=8'd244;
		data_a[15588]<=8'd244;
		data_a[15589]<=8'd244;
		data_a[15590]<=8'd243;
		data_a[15591]<=8'd244;
		data_a[15592]<=8'd246;
		data_a[15593]<=8'd248;
		data_a[15594]<=8'd246;
		data_a[15595]<=8'd246;
		data_a[15596]<=8'd247;
		data_a[15597]<=8'd247;
		data_a[15598]<=8'd247;
		data_a[15599]<=8'd247;
		data_a[15600]<=8'd255;
		data_a[15601]<=8'd83;
		data_a[15602]<=8'd84;
		data_a[15603]<=8'd84;
		data_a[15604]<=8'd81;
		data_a[15605]<=8'd80;
		data_a[15606]<=8'd79;
		data_a[15607]<=8'd70;
		data_a[15608]<=8'd74;
		data_a[15609]<=8'd65;
		data_a[15610]<=8'd62;
		data_a[15611]<=8'd75;
		data_a[15612]<=8'd75;
		data_a[15613]<=8'd67;
		data_a[15614]<=8'd73;
		data_a[15615]<=8'd72;
		data_a[15616]<=8'd70;
		data_a[15617]<=8'd62;
		data_a[15618]<=8'd55;
		data_a[15619]<=8'd59;
		data_a[15620]<=8'd53;
		data_a[15621]<=8'd156;
		data_a[15622]<=8'd137;
		data_a[15623]<=8'd145;
		data_a[15624]<=8'd141;
		data_a[15625]<=8'd67;
		data_a[15626]<=8'd57;
		data_a[15627]<=8'd57;
		data_a[15628]<=8'd109;
		data_a[15629]<=8'd137;
		data_a[15630]<=8'd131;
		data_a[15631]<=8'd131;
		data_a[15632]<=8'd130;
		data_a[15633]<=8'd121;
		data_a[15634]<=8'd120;
		data_a[15635]<=8'd105;
		data_a[15636]<=8'd97;
		data_a[15637]<=8'd85;
		data_a[15638]<=8'd106;
		data_a[15639]<=8'd116;
		data_a[15640]<=8'd117;
		data_a[15641]<=8'd114;
		data_a[15642]<=8'd104;
		data_a[15643]<=8'd107;
		data_a[15644]<=8'd111;
		data_a[15645]<=8'd119;
		data_a[15646]<=8'd124;
		data_a[15647]<=8'd110;
		data_a[15648]<=8'd111;
		data_a[15649]<=8'd119;
		data_a[15650]<=8'd113;
		data_a[15651]<=8'd120;
		data_a[15652]<=8'd115;
		data_a[15653]<=8'd90;
		data_a[15654]<=8'd90;
		data_a[15655]<=8'd100;
		data_a[15656]<=8'd114;
		data_a[15657]<=8'd115;
		data_a[15658]<=8'd114;
		data_a[15659]<=8'd127;
		data_a[15660]<=8'd123;
		data_a[15661]<=8'd144;
		data_a[15662]<=8'd153;
		data_a[15663]<=8'd149;
		data_a[15664]<=8'd104;
		data_a[15665]<=8'd147;
		data_a[15666]<=8'd190;
		data_a[15667]<=8'd184;
		data_a[15668]<=8'd218;
		data_a[15669]<=8'd221;
		data_a[15670]<=8'd225;
		data_a[15671]<=8'd224;
		data_a[15672]<=8'd224;
		data_a[15673]<=8'd230;
		data_a[15674]<=8'd223;
		data_a[15675]<=8'd229;
		data_a[15676]<=8'd223;
		data_a[15677]<=8'd239;
		data_a[15678]<=8'd235;
		data_a[15679]<=8'd237;
		data_a[15680]<=8'd234;
		data_a[15681]<=8'd239;
		data_a[15682]<=8'd228;
		data_a[15683]<=8'd238;
		data_a[15684]<=8'd142;
		data_a[15685]<=8'd82;
		data_a[15686]<=8'd74;
		data_a[15687]<=8'd104;
		data_a[15688]<=8'd122;
		data_a[15689]<=8'd129;
		data_a[15690]<=8'd142;
		data_a[15691]<=8'd141;
		data_a[15692]<=8'd116;
		data_a[15693]<=8'd69;
		data_a[15694]<=8'd69;
		data_a[15695]<=8'd68;
		data_a[15696]<=8'd61;
		data_a[15697]<=8'd62;
		data_a[15698]<=8'd59;
		data_a[15699]<=8'd66;
		data_a[15700]<=8'd66;
		data_a[15701]<=8'd82;
		data_a[15702]<=8'd90;
		data_a[15703]<=8'd97;
		data_a[15704]<=8'd115;
		data_a[15705]<=8'd126;
		data_a[15706]<=8'd122;
		data_a[15707]<=8'd125;
		data_a[15708]<=8'd117;
		data_a[15709]<=8'd116;
		data_a[15710]<=8'd124;
		data_a[15711]<=8'd126;
		data_a[15712]<=8'd137;
		data_a[15713]<=8'd134;
		data_a[15714]<=8'd139;
		data_a[15715]<=8'd132;
		data_a[15716]<=8'd135;
		data_a[15717]<=8'd127;
		data_a[15718]<=8'd117;
		data_a[15719]<=8'd106;
		data_a[15720]<=8'd101;
		data_a[15721]<=8'd94;
		data_a[15722]<=8'd107;
		data_a[15723]<=8'd95;
		data_a[15724]<=8'd72;
		data_a[15725]<=8'd65;
		data_a[15726]<=8'd64;
		data_a[15727]<=8'd65;
		data_a[15728]<=8'd59;
		data_a[15729]<=8'd73;
		data_a[15730]<=8'd68;
		data_a[15731]<=8'd83;
		data_a[15732]<=8'd131;
		data_a[15733]<=8'd183;
		data_a[15734]<=8'd237;
		data_a[15735]<=8'd245;
		data_a[15736]<=8'd244;
		data_a[15737]<=8'd243;
		data_a[15738]<=8'd244;
		data_a[15739]<=8'd243;
		data_a[15740]<=8'd246;
		data_a[15741]<=8'd247;
		data_a[15742]<=8'd243;
		data_a[15743]<=8'd245;
		data_a[15744]<=8'd247;
		data_a[15745]<=8'd249;
		data_a[15746]<=8'd248;
		data_a[15747]<=8'd246;
		data_a[15748]<=8'd248;
		data_a[15749]<=8'd248;
		data_a[15750]<=8'd255;
		data_a[15751]<=8'd85;
		data_a[15752]<=8'd86;
		data_a[15753]<=8'd83;
		data_a[15754]<=8'd79;
		data_a[15755]<=8'd78;
		data_a[15756]<=8'd79;
		data_a[15757]<=8'd71;
		data_a[15758]<=8'd132;
		data_a[15759]<=8'd65;
		data_a[15760]<=8'd69;
		data_a[15761]<=8'd74;
		data_a[15762]<=8'd75;
		data_a[15763]<=8'd73;
		data_a[15764]<=8'd72;
		data_a[15765]<=8'd69;
		data_a[15766]<=8'd64;
		data_a[15767]<=8'd68;
		data_a[15768]<=8'd55;
		data_a[15769]<=8'd62;
		data_a[15770]<=8'd39;
		data_a[15771]<=8'd147;
		data_a[15772]<=8'd141;
		data_a[15773]<=8'd142;
		data_a[15774]<=8'd150;
		data_a[15775]<=8'd110;
		data_a[15776]<=8'd82;
		data_a[15777]<=8'd53;
		data_a[15778]<=8'd103;
		data_a[15779]<=8'd135;
		data_a[15780]<=8'd126;
		data_a[15781]<=8'd123;
		data_a[15782]<=8'd124;
		data_a[15783]<=8'd125;
		data_a[15784]<=8'd121;
		data_a[15785]<=8'd106;
		data_a[15786]<=8'd91;
		data_a[15787]<=8'd88;
		data_a[15788]<=8'd104;
		data_a[15789]<=8'd110;
		data_a[15790]<=8'd120;
		data_a[15791]<=8'd117;
		data_a[15792]<=8'd100;
		data_a[15793]<=8'd85;
		data_a[15794]<=8'd82;
		data_a[15795]<=8'd102;
		data_a[15796]<=8'd108;
		data_a[15797]<=8'd101;
		data_a[15798]<=8'd109;
		data_a[15799]<=8'd109;
		data_a[15800]<=8'd86;
		data_a[15801]<=8'd98;
		data_a[15802]<=8'd96;
		data_a[15803]<=8'd98;
		data_a[15804]<=8'd90;
		data_a[15805]<=8'd97;
		data_a[15806]<=8'd104;
		data_a[15807]<=8'd109;
		data_a[15808]<=8'd116;
		data_a[15809]<=8'd119;
		data_a[15810]<=8'd125;
		data_a[15811]<=8'd147;
		data_a[15812]<=8'd137;
		data_a[15813]<=8'd148;
		data_a[15814]<=8'd111;
		data_a[15815]<=8'd183;
		data_a[15816]<=8'd124;
		data_a[15817]<=8'd198;
		data_a[15818]<=8'd226;
		data_a[15819]<=8'd222;
		data_a[15820]<=8'd228;
		data_a[15821]<=8'd230;
		data_a[15822]<=8'd227;
		data_a[15823]<=8'd230;
		data_a[15824]<=8'd226;
		data_a[15825]<=8'd228;
		data_a[15826]<=8'd226;
		data_a[15827]<=8'd238;
		data_a[15828]<=8'd238;
		data_a[15829]<=8'd238;
		data_a[15830]<=8'd233;
		data_a[15831]<=8'd237;
		data_a[15832]<=8'd240;
		data_a[15833]<=8'd229;
		data_a[15834]<=8'd110;
		data_a[15835]<=8'd77;
		data_a[15836]<=8'd71;
		data_a[15837]<=8'd101;
		data_a[15838]<=8'd113;
		data_a[15839]<=8'd130;
		data_a[15840]<=8'd135;
		data_a[15841]<=8'd137;
		data_a[15842]<=8'd125;
		data_a[15843]<=8'd81;
		data_a[15844]<=8'd70;
		data_a[15845]<=8'd62;
		data_a[15846]<=8'd59;
		data_a[15847]<=8'd55;
		data_a[15848]<=8'd63;
		data_a[15849]<=8'd72;
		data_a[15850]<=8'd89;
		data_a[15851]<=8'd98;
		data_a[15852]<=8'd113;
		data_a[15853]<=8'd119;
		data_a[15854]<=8'd124;
		data_a[15855]<=8'd121;
		data_a[15856]<=8'd119;
		data_a[15857]<=8'd111;
		data_a[15858]<=8'd115;
		data_a[15859]<=8'd118;
		data_a[15860]<=8'd127;
		data_a[15861]<=8'd129;
		data_a[15862]<=8'd128;
		data_a[15863]<=8'd128;
		data_a[15864]<=8'd128;
		data_a[15865]<=8'd133;
		data_a[15866]<=8'd133;
		data_a[15867]<=8'd136;
		data_a[15868]<=8'd123;
		data_a[15869]<=8'd117;
		data_a[15870]<=8'd105;
		data_a[15871]<=8'd96;
		data_a[15872]<=8'd100;
		data_a[15873]<=8'd89;
		data_a[15874]<=8'd72;
		data_a[15875]<=8'd62;
		data_a[15876]<=8'd64;
		data_a[15877]<=8'd58;
		data_a[15878]<=8'd65;
		data_a[15879]<=8'd65;
		data_a[15880]<=8'd69;
		data_a[15881]<=8'd79;
		data_a[15882]<=8'd117;
		data_a[15883]<=8'd209;
		data_a[15884]<=8'd247;
		data_a[15885]<=8'd241;
		data_a[15886]<=8'd244;
		data_a[15887]<=8'd244;
		data_a[15888]<=8'd246;
		data_a[15889]<=8'd244;
		data_a[15890]<=8'd246;
		data_a[15891]<=8'd247;
		data_a[15892]<=8'd244;
		data_a[15893]<=8'd246;
		data_a[15894]<=8'd245;
		data_a[15895]<=8'd247;
		data_a[15896]<=8'd247;
		data_a[15897]<=8'd246;
		data_a[15898]<=8'd247;
		data_a[15899]<=8'd247;
		data_a[15900]<=8'd254;
		data_a[15901]<=8'd83;
		data_a[15902]<=8'd86;
		data_a[15903]<=8'd85;
		data_a[15904]<=8'd82;
		data_a[15905]<=8'd83;
		data_a[15906]<=8'd86;
		data_a[15907]<=8'd79;
		data_a[15908]<=8'd140;
		data_a[15909]<=8'd92;
		data_a[15910]<=8'd67;
		data_a[15911]<=8'd72;
		data_a[15912]<=8'd68;
		data_a[15913]<=8'd69;
		data_a[15914]<=8'd69;
		data_a[15915]<=8'd71;
		data_a[15916]<=8'd68;
		data_a[15917]<=8'd65;
		data_a[15918]<=8'd49;
		data_a[15919]<=8'd84;
		data_a[15920]<=8'd54;
		data_a[15921]<=8'd147;
		data_a[15922]<=8'd145;
		data_a[15923]<=8'd146;
		data_a[15924]<=8'd146;
		data_a[15925]<=8'd143;
		data_a[15926]<=8'd98;
		data_a[15927]<=8'd68;
		data_a[15928]<=8'd102;
		data_a[15929]<=8'd132;
		data_a[15930]<=8'd119;
		data_a[15931]<=8'd123;
		data_a[15932]<=8'd117;
		data_a[15933]<=8'd120;
		data_a[15934]<=8'd113;
		data_a[15935]<=8'd94;
		data_a[15936]<=8'd85;
		data_a[15937]<=8'd91;
		data_a[15938]<=8'd106;
		data_a[15939]<=8'd107;
		data_a[15940]<=8'd115;
		data_a[15941]<=8'd105;
		data_a[15942]<=8'd102;
		data_a[15943]<=8'd100;
		data_a[15944]<=8'd82;
		data_a[15945]<=8'd93;
		data_a[15946]<=8'd96;
		data_a[15947]<=8'd93;
		data_a[15948]<=8'd97;
		data_a[15949]<=8'd92;
		data_a[15950]<=8'd88;
		data_a[15951]<=8'd81;
		data_a[15952]<=8'd101;
		data_a[15953]<=8'd97;
		data_a[15954]<=8'd96;
		data_a[15955]<=8'd90;
		data_a[15956]<=8'd104;
		data_a[15957]<=8'd105;
		data_a[15958]<=8'd118;
		data_a[15959]<=8'd115;
		data_a[15960]<=8'd125;
		data_a[15961]<=8'd135;
		data_a[15962]<=8'd150;
		data_a[15963]<=8'd125;
		data_a[15964]<=8'd137;
		data_a[15965]<=8'd168;
		data_a[15966]<=8'd89;
		data_a[15967]<=8'd227;
		data_a[15968]<=8'd223;
		data_a[15969]<=8'd224;
		data_a[15970]<=8'd226;
		data_a[15971]<=8'd224;
		data_a[15972]<=8'd227;
		data_a[15973]<=8'd230;
		data_a[15974]<=8'd229;
		data_a[15975]<=8'd228;
		data_a[15976]<=8'd229;
		data_a[15977]<=8'd236;
		data_a[15978]<=8'd239;
		data_a[15979]<=8'd238;
		data_a[15980]<=8'd239;
		data_a[15981]<=8'd235;
		data_a[15982]<=8'd235;
		data_a[15983]<=8'd235;
		data_a[15984]<=8'd209;
		data_a[15985]<=8'd83;
		data_a[15986]<=8'd76;
		data_a[15987]<=8'd86;
		data_a[15988]<=8'd96;
		data_a[15989]<=8'd119;
		data_a[15990]<=8'd125;
		data_a[15991]<=8'd134;
		data_a[15992]<=8'd138;
		data_a[15993]<=8'd65;
		data_a[15994]<=8'd66;
		data_a[15995]<=8'd63;
		data_a[15996]<=8'd62;
		data_a[15997]<=8'd63;
		data_a[15998]<=8'd64;
		data_a[15999]<=8'd79;
		data_a[16000]<=8'd87;
		data_a[16001]<=8'd100;
		data_a[16002]<=8'd103;
		data_a[16003]<=8'd108;
		data_a[16004]<=8'd112;
		data_a[16005]<=8'd111;
		data_a[16006]<=8'd121;
		data_a[16007]<=8'd119;
		data_a[16008]<=8'd127;
		data_a[16009]<=8'd129;
		data_a[16010]<=8'd124;
		data_a[16011]<=8'd121;
		data_a[16012]<=8'd119;
		data_a[16013]<=8'd114;
		data_a[16014]<=8'd124;
		data_a[16015]<=8'd122;
		data_a[16016]<=8'd136;
		data_a[16017]<=8'd131;
		data_a[16018]<=8'd129;
		data_a[16019]<=8'd121;
		data_a[16020]<=8'd104;
		data_a[16021]<=8'd100;
		data_a[16022]<=8'd96;
		data_a[16023]<=8'd89;
		data_a[16024]<=8'd67;
		data_a[16025]<=8'd59;
		data_a[16026]<=8'd64;
		data_a[16027]<=8'd61;
		data_a[16028]<=8'd66;
		data_a[16029]<=8'd61;
		data_a[16030]<=8'd76;
		data_a[16031]<=8'd94;
		data_a[16032]<=8'd128;
		data_a[16033]<=8'd178;
		data_a[16034]<=8'd246;
		data_a[16035]<=8'd243;
		data_a[16036]<=8'd245;
		data_a[16037]<=8'd245;
		data_a[16038]<=8'd247;
		data_a[16039]<=8'd246;
		data_a[16040]<=8'd247;
		data_a[16041]<=8'd248;
		data_a[16042]<=8'd245;
		data_a[16043]<=8'd248;
		data_a[16044]<=8'd245;
		data_a[16045]<=8'd248;
		data_a[16046]<=8'd247;
		data_a[16047]<=8'd246;
		data_a[16048]<=8'd248;
		data_a[16049]<=8'd248;
		data_a[16050]<=8'd254;
		data_a[16051]<=8'd83;
		data_a[16052]<=8'd86;
		data_a[16053]<=8'd85;
		data_a[16054]<=8'd82;
		data_a[16055]<=8'd81;
		data_a[16056]<=8'd80;
		data_a[16057]<=8'd69;
		data_a[16058]<=8'd109;
		data_a[16059]<=8'd104;
		data_a[16060]<=8'd61;
		data_a[16061]<=8'd72;
		data_a[16062]<=8'd75;
		data_a[16063]<=8'd73;
		data_a[16064]<=8'd75;
		data_a[16065]<=8'd75;
		data_a[16066]<=8'd71;
		data_a[16067]<=8'd68;
		data_a[16068]<=8'd49;
		data_a[16069]<=8'd81;
		data_a[16070]<=8'd56;
		data_a[16071]<=8'd149;
		data_a[16072]<=8'd152;
		data_a[16073]<=8'd147;
		data_a[16074]<=8'd149;
		data_a[16075]<=8'd155;
		data_a[16076]<=8'd93;
		data_a[16077]<=8'd69;
		data_a[16078]<=8'd94;
		data_a[16079]<=8'd122;
		data_a[16080]<=8'd126;
		data_a[16081]<=8'd124;
		data_a[16082]<=8'd119;
		data_a[16083]<=8'd115;
		data_a[16084]<=8'd107;
		data_a[16085]<=8'd86;
		data_a[16086]<=8'd91;
		data_a[16087]<=8'd94;
		data_a[16088]<=8'd111;
		data_a[16089]<=8'd107;
		data_a[16090]<=8'd109;
		data_a[16091]<=8'd106;
		data_a[16092]<=8'd86;
		data_a[16093]<=8'd77;
		data_a[16094]<=8'd82;
		data_a[16095]<=8'd90;
		data_a[16096]<=8'd85;
		data_a[16097]<=8'd83;
		data_a[16098]<=8'd78;
		data_a[16099]<=8'd77;
		data_a[16100]<=8'd79;
		data_a[16101]<=8'd77;
		data_a[16102]<=8'd95;
		data_a[16103]<=8'd101;
		data_a[16104]<=8'd97;
		data_a[16105]<=8'd94;
		data_a[16106]<=8'd96;
		data_a[16107]<=8'd97;
		data_a[16108]<=8'd102;
		data_a[16109]<=8'd114;
		data_a[16110]<=8'd125;
		data_a[16111]<=8'd143;
		data_a[16112]<=8'd134;
		data_a[16113]<=8'd111;
		data_a[16114]<=8'd161;
		data_a[16115]<=8'd123;
		data_a[16116]<=8'd97;
		data_a[16117]<=8'd224;
		data_a[16118]<=8'd226;
		data_a[16119]<=8'd230;
		data_a[16120]<=8'd226;
		data_a[16121]<=8'd226;
		data_a[16122]<=8'd227;
		data_a[16123]<=8'd230;
		data_a[16124]<=8'd230;
		data_a[16125]<=8'd231;
		data_a[16126]<=8'd231;
		data_a[16127]<=8'd237;
		data_a[16128]<=8'd239;
		data_a[16129]<=8'd238;
		data_a[16130]<=8'd236;
		data_a[16131]<=8'd236;
		data_a[16132]<=8'd235;
		data_a[16133]<=8'd235;
		data_a[16134]<=8'd231;
		data_a[16135]<=8'd120;
		data_a[16136]<=8'd77;
		data_a[16137]<=8'd77;
		data_a[16138]<=8'd88;
		data_a[16139]<=8'd106;
		data_a[16140]<=8'd122;
		data_a[16141]<=8'd131;
		data_a[16142]<=8'd133;
		data_a[16143]<=8'd96;
		data_a[16144]<=8'd63;
		data_a[16145]<=8'd67;
		data_a[16146]<=8'd74;
		data_a[16147]<=8'd75;
		data_a[16148]<=8'd79;
		data_a[16149]<=8'd74;
		data_a[16150]<=8'd90;
		data_a[16151]<=8'd99;
		data_a[16152]<=8'd110;
		data_a[16153]<=8'd108;
		data_a[16154]<=8'd117;
		data_a[16155]<=8'd118;
		data_a[16156]<=8'd122;
		data_a[16157]<=8'd121;
		data_a[16158]<=8'd115;
		data_a[16159]<=8'd117;
		data_a[16160]<=8'd106;
		data_a[16161]<=8'd107;
		data_a[16162]<=8'd109;
		data_a[16163]<=8'd110;
		data_a[16164]<=8'd118;
		data_a[16165]<=8'd123;
		data_a[16166]<=8'd129;
		data_a[16167]<=8'd131;
		data_a[16168]<=8'd126;
		data_a[16169]<=8'd123;
		data_a[16170]<=8'd108;
		data_a[16171]<=8'd98;
		data_a[16172]<=8'd87;
		data_a[16173]<=8'd86;
		data_a[16174]<=8'd67;
		data_a[16175]<=8'd68;
		data_a[16176]<=8'd64;
		data_a[16177]<=8'd61;
		data_a[16178]<=8'd65;
		data_a[16179]<=8'd74;
		data_a[16180]<=8'd78;
		data_a[16181]<=8'd78;
		data_a[16182]<=8'd116;
		data_a[16183]<=8'd115;
		data_a[16184]<=8'd248;
		data_a[16185]<=8'd247;
		data_a[16186]<=8'd245;
		data_a[16187]<=8'd246;
		data_a[16188]<=8'd248;
		data_a[16189]<=8'd246;
		data_a[16190]<=8'd247;
		data_a[16191]<=8'd248;
		data_a[16192]<=8'd245;
		data_a[16193]<=8'd249;
		data_a[16194]<=8'd247;
		data_a[16195]<=8'd249;
		data_a[16196]<=8'd248;
		data_a[16197]<=8'd246;
		data_a[16198]<=8'd248;
		data_a[16199]<=8'd250;
		data_a[16200]<=8'd255;
		data_a[16201]<=8'd84;
		data_a[16202]<=8'd84;
		data_a[16203]<=8'd84;
		data_a[16204]<=8'd83;
		data_a[16205]<=8'd82;
		data_a[16206]<=8'd76;
		data_a[16207]<=8'd62;
		data_a[16208]<=8'd78;
		data_a[16209]<=8'd69;
		data_a[16210]<=8'd65;
		data_a[16211]<=8'd71;
		data_a[16212]<=8'd73;
		data_a[16213]<=8'd68;
		data_a[16214]<=8'd72;
		data_a[16215]<=8'd73;
		data_a[16216]<=8'd71;
		data_a[16217]<=8'd68;
		data_a[16218]<=8'd53;
		data_a[16219]<=8'd69;
		data_a[16220]<=8'd51;
		data_a[16221]<=8'd143;
		data_a[16222]<=8'd151;
		data_a[16223]<=8'd147;
		data_a[16224]<=8'd152;
		data_a[16225]<=8'd143;
		data_a[16226]<=8'd134;
		data_a[16227]<=8'd77;
		data_a[16228]<=8'd78;
		data_a[16229]<=8'd123;
		data_a[16230]<=8'd116;
		data_a[16231]<=8'd126;
		data_a[16232]<=8'd120;
		data_a[16233]<=8'd112;
		data_a[16234]<=8'd103;
		data_a[16235]<=8'd88;
		data_a[16236]<=8'd96;
		data_a[16237]<=8'd93;
		data_a[16238]<=8'd107;
		data_a[16239]<=8'd106;
		data_a[16240]<=8'd105;
		data_a[16241]<=8'd103;
		data_a[16242]<=8'd85;
		data_a[16243]<=8'd74;
		data_a[16244]<=8'd67;
		data_a[16245]<=8'd59;
		data_a[16246]<=8'd72;
		data_a[16247]<=8'd71;
		data_a[16248]<=8'd72;
		data_a[16249]<=8'd65;
		data_a[16250]<=8'd74;
		data_a[16251]<=8'd73;
		data_a[16252]<=8'd98;
		data_a[16253]<=8'd101;
		data_a[16254]<=8'd95;
		data_a[16255]<=8'd88;
		data_a[16256]<=8'd87;
		data_a[16257]<=8'd102;
		data_a[16258]<=8'd107;
		data_a[16259]<=8'd113;
		data_a[16260]<=8'd118;
		data_a[16261]<=8'd138;
		data_a[16262]<=8'd137;
		data_a[16263]<=8'd96;
		data_a[16264]<=8'd132;
		data_a[16265]<=8'd162;
		data_a[16266]<=8'd192;
		data_a[16267]<=8'd226;
		data_a[16268]<=8'd224;
		data_a[16269]<=8'd223;
		data_a[16270]<=8'd229;
		data_a[16271]<=8'd234;
		data_a[16272]<=8'd228;
		data_a[16273]<=8'd232;
		data_a[16274]<=8'd230;
		data_a[16275]<=8'd233;
		data_a[16276]<=8'd231;
		data_a[16277]<=8'd239;
		data_a[16278]<=8'd239;
		data_a[16279]<=8'd240;
		data_a[16280]<=8'd237;
		data_a[16281]<=8'd235;
		data_a[16282]<=8'd246;
		data_a[16283]<=8'd239;
		data_a[16284]<=8'd234;
		data_a[16285]<=8'd123;
		data_a[16286]<=8'd69;
		data_a[16287]<=8'd86;
		data_a[16288]<=8'd82;
		data_a[16289]<=8'd82;
		data_a[16290]<=8'd110;
		data_a[16291]<=8'd126;
		data_a[16292]<=8'd140;
		data_a[16293]<=8'd104;
		data_a[16294]<=8'd71;
		data_a[16295]<=8'd66;
		data_a[16296]<=8'd69;
		data_a[16297]<=8'd83;
		data_a[16298]<=8'd99;
		data_a[16299]<=8'd99;
		data_a[16300]<=8'd115;
		data_a[16301]<=8'd118;
		data_a[16302]<=8'd121;
		data_a[16303]<=8'd114;
		data_a[16304]<=8'd123;
		data_a[16305]<=8'd118;
		data_a[16306]<=8'd107;
		data_a[16307]<=8'd100;
		data_a[16308]<=8'd88;
		data_a[16309]<=8'd88;
		data_a[16310]<=8'd90;
		data_a[16311]<=8'd96;
		data_a[16312]<=8'd103;
		data_a[16313]<=8'd109;
		data_a[16314]<=8'd120;
		data_a[16315]<=8'd125;
		data_a[16316]<=8'd129;
		data_a[16317]<=8'd131;
		data_a[16318]<=8'd128;
		data_a[16319]<=8'd126;
		data_a[16320]<=8'd107;
		data_a[16321]<=8'd95;
		data_a[16322]<=8'd91;
		data_a[16323]<=8'd80;
		data_a[16324]<=8'd66;
		data_a[16325]<=8'd66;
		data_a[16326]<=8'd61;
		data_a[16327]<=8'd62;
		data_a[16328]<=8'd60;
		data_a[16329]<=8'd76;
		data_a[16330]<=8'd77;
		data_a[16331]<=8'd89;
		data_a[16332]<=8'd85;
		data_a[16333]<=8'd167;
		data_a[16334]<=8'd239;
		data_a[16335]<=8'd246;
		data_a[16336]<=8'd245;
		data_a[16337]<=8'd246;
		data_a[16338]<=8'd248;
		data_a[16339]<=8'd246;
		data_a[16340]<=8'd247;
		data_a[16341]<=8'd248;
		data_a[16342]<=8'd245;
		data_a[16343]<=8'd248;
		data_a[16344]<=8'd247;
		data_a[16345]<=8'd248;
		data_a[16346]<=8'd247;
		data_a[16347]<=8'd245;
		data_a[16348]<=8'd247;
		data_a[16349]<=8'd248;
		data_a[16350]<=8'd255;
		data_a[16351]<=8'd82;
		data_a[16352]<=8'd81;
		data_a[16353]<=8'd82;
		data_a[16354]<=8'd84;
		data_a[16355]<=8'd86;
		data_a[16356]<=8'd80;
		data_a[16357]<=8'd64;
		data_a[16358]<=8'd66;
		data_a[16359]<=8'd58;
		data_a[16360]<=8'd72;
		data_a[16361]<=8'd79;
		data_a[16362]<=8'd71;
		data_a[16363]<=8'd72;
		data_a[16364]<=8'd73;
		data_a[16365]<=8'd74;
		data_a[16366]<=8'd71;
		data_a[16367]<=8'd65;
		data_a[16368]<=8'd51;
		data_a[16369]<=8'd68;
		data_a[16370]<=8'd51;
		data_a[16371]<=8'd145;
		data_a[16372]<=8'd151;
		data_a[16373]<=8'd148;
		data_a[16374]<=8'd145;
		data_a[16375]<=8'd155;
		data_a[16376]<=8'd155;
		data_a[16377]<=8'd131;
		data_a[16378]<=8'd94;
		data_a[16379]<=8'd121;
		data_a[16380]<=8'd119;
		data_a[16381]<=8'd119;
		data_a[16382]<=8'd116;
		data_a[16383]<=8'd111;
		data_a[16384]<=8'd99;
		data_a[16385]<=8'd90;
		data_a[16386]<=8'd91;
		data_a[16387]<=8'd92;
		data_a[16388]<=8'd105;
		data_a[16389]<=8'd113;
		data_a[16390]<=8'd119;
		data_a[16391]<=8'd124;
		data_a[16392]<=8'd105;
		data_a[16393]<=8'd107;
		data_a[16394]<=8'd117;
		data_a[16395]<=8'd80;
		data_a[16396]<=8'd65;
		data_a[16397]<=8'd56;
		data_a[16398]<=8'd62;
		data_a[16399]<=8'd58;
		data_a[16400]<=8'd63;
		data_a[16401]<=8'd74;
		data_a[16402]<=8'd91;
		data_a[16403]<=8'd99;
		data_a[16404]<=8'd89;
		data_a[16405]<=8'd85;
		data_a[16406]<=8'd82;
		data_a[16407]<=8'd91;
		data_a[16408]<=8'd101;
		data_a[16409]<=8'd110;
		data_a[16410]<=8'd130;
		data_a[16411]<=8'd132;
		data_a[16412]<=8'd145;
		data_a[16413]<=8'd78;
		data_a[16414]<=8'd201;
		data_a[16415]<=8'd204;
		data_a[16416]<=8'd216;
		data_a[16417]<=8'd222;
		data_a[16418]<=8'd231;
		data_a[16419]<=8'd230;
		data_a[16420]<=8'd229;
		data_a[16421]<=8'd229;
		data_a[16422]<=8'd230;
		data_a[16423]<=8'd232;
		data_a[16424]<=8'd228;
		data_a[16425]<=8'd231;
		data_a[16426]<=8'd230;
		data_a[16427]<=8'd240;
		data_a[16428]<=8'd240;
		data_a[16429]<=8'd241;
		data_a[16430]<=8'd240;
		data_a[16431]<=8'd239;
		data_a[16432]<=8'd231;
		data_a[16433]<=8'd238;
		data_a[16434]<=8'd215;
		data_a[16435]<=8'd124;
		data_a[16436]<=8'd84;
		data_a[16437]<=8'd77;
		data_a[16438]<=8'd77;
		data_a[16439]<=8'd80;
		data_a[16440]<=8'd116;
		data_a[16441]<=8'd122;
		data_a[16442]<=8'd126;
		data_a[16443]<=8'd138;
		data_a[16444]<=8'd82;
		data_a[16445]<=8'd65;
		data_a[16446]<=8'd74;
		data_a[16447]<=8'd92;
		data_a[16448]<=8'd101;
		data_a[16449]<=8'd111;
		data_a[16450]<=8'd114;
		data_a[16451]<=8'd122;
		data_a[16452]<=8'd118;
		data_a[16453]<=8'd120;
		data_a[16454]<=8'd108;
		data_a[16455]<=8'd96;
		data_a[16456]<=8'd86;
		data_a[16457]<=8'd77;
		data_a[16458]<=8'd77;
		data_a[16459]<=8'd73;
		data_a[16460]<=8'd82;
		data_a[16461]<=8'd88;
		data_a[16462]<=8'd100;
		data_a[16463]<=8'd107;
		data_a[16464]<=8'd126;
		data_a[16465]<=8'd123;
		data_a[16466]<=8'd134;
		data_a[16467]<=8'd129;
		data_a[16468]<=8'd131;
		data_a[16469]<=8'd125;
		data_a[16470]<=8'd104;
		data_a[16471]<=8'd93;
		data_a[16472]<=8'd102;
		data_a[16473]<=8'd76;
		data_a[16474]<=8'd66;
		data_a[16475]<=8'd54;
		data_a[16476]<=8'd60;
		data_a[16477]<=8'd65;
		data_a[16478]<=8'd65;
		data_a[16479]<=8'd65;
		data_a[16480]<=8'd74;
		data_a[16481]<=8'd77;
		data_a[16482]<=8'd84;
		data_a[16483]<=8'd134;
		data_a[16484]<=8'd251;
		data_a[16485]<=8'd240;
		data_a[16486]<=8'd245;
		data_a[16487]<=8'd245;
		data_a[16488]<=8'd247;
		data_a[16489]<=8'd246;
		data_a[16490]<=8'd247;
		data_a[16491]<=8'd248;
		data_a[16492]<=8'd245;
		data_a[16493]<=8'd248;
		data_a[16494]<=8'd245;
		data_a[16495]<=8'd248;
		data_a[16496]<=8'd247;
		data_a[16497]<=8'd246;
		data_a[16498]<=8'd247;
		data_a[16499]<=8'd247;
		data_a[16500]<=8'd255;
		data_a[16501]<=8'd82;
		data_a[16502]<=8'd81;
		data_a[16503]<=8'd79;
		data_a[16504]<=8'd79;
		data_a[16505]<=8'd79;
		data_a[16506]<=8'd72;
		data_a[16507]<=8'd56;
		data_a[16508]<=8'd59;
		data_a[16509]<=8'd62;
		data_a[16510]<=8'd63;
		data_a[16511]<=8'd73;
		data_a[16512]<=8'd71;
		data_a[16513]<=8'd75;
		data_a[16514]<=8'd71;
		data_a[16515]<=8'd67;
		data_a[16516]<=8'd70;
		data_a[16517]<=8'd69;
		data_a[16518]<=8'd50;
		data_a[16519]<=8'd75;
		data_a[16520]<=8'd44;
		data_a[16521]<=8'd151;
		data_a[16522]<=8'd158;
		data_a[16523]<=8'd150;
		data_a[16524]<=8'd158;
		data_a[16525]<=8'd161;
		data_a[16526]<=8'd153;
		data_a[16527]<=8'd162;
		data_a[16528]<=8'd118;
		data_a[16529]<=8'd126;
		data_a[16530]<=8'd118;
		data_a[16531]<=8'd117;
		data_a[16532]<=8'd115;
		data_a[16533]<=8'd114;
		data_a[16534]<=8'd101;
		data_a[16535]<=8'd89;
		data_a[16536]<=8'd89;
		data_a[16537]<=8'd91;
		data_a[16538]<=8'd102;
		data_a[16539]<=8'd108;
		data_a[16540]<=8'd103;
		data_a[16541]<=8'd107;
		data_a[16542]<=8'd99;
		data_a[16543]<=8'd97;
		data_a[16544]<=8'd101;
		data_a[16545]<=8'd96;
		data_a[16546]<=8'd102;
		data_a[16547]<=8'd87;
		data_a[16548]<=8'd92;
		data_a[16549]<=8'd81;
		data_a[16550]<=8'd90;
		data_a[16551]<=8'd81;
		data_a[16552]<=8'd99;
		data_a[16553]<=8'd86;
		data_a[16554]<=8'd87;
		data_a[16555]<=8'd79;
		data_a[16556]<=8'd85;
		data_a[16557]<=8'd93;
		data_a[16558]<=8'd101;
		data_a[16559]<=8'd113;
		data_a[16560]<=8'd127;
		data_a[16561]<=8'd130;
		data_a[16562]<=8'd135;
		data_a[16563]<=8'd157;
		data_a[16564]<=8'd230;
		data_a[16565]<=8'd215;
		data_a[16566]<=8'd223;
		data_a[16567]<=8'd228;
		data_a[16568]<=8'd225;
		data_a[16569]<=8'd230;
		data_a[16570]<=8'd229;
		data_a[16571]<=8'd227;
		data_a[16572]<=8'd230;
		data_a[16573]<=8'd230;
		data_a[16574]<=8'd230;
		data_a[16575]<=8'd231;
		data_a[16576]<=8'd234;
		data_a[16577]<=8'd240;
		data_a[16578]<=8'd242;
		data_a[16579]<=8'd241;
		data_a[16580]<=8'd238;
		data_a[16581]<=8'd244;
		data_a[16582]<=8'd237;
		data_a[16583]<=8'd234;
		data_a[16584]<=8'd234;
		data_a[16585]<=8'd169;
		data_a[16586]<=8'd77;
		data_a[16587]<=8'd79;
		data_a[16588]<=8'd79;
		data_a[16589]<=8'd72;
		data_a[16590]<=8'd92;
		data_a[16591]<=8'd106;
		data_a[16592]<=8'd130;
		data_a[16593]<=8'd130;
		data_a[16594]<=8'd99;
		data_a[16595]<=8'd66;
		data_a[16596]<=8'd78;
		data_a[16597]<=8'd96;
		data_a[16598]<=8'd112;
		data_a[16599]<=8'd112;
		data_a[16600]<=8'd122;
		data_a[16601]<=8'd116;
		data_a[16602]<=8'd111;
		data_a[16603]<=8'd106;
		data_a[16604]<=8'd97;
		data_a[16605]<=8'd80;
		data_a[16606]<=8'd74;
		data_a[16607]<=8'd66;
		data_a[16608]<=8'd69;
		data_a[16609]<=8'd68;
		data_a[16610]<=8'd75;
		data_a[16611]<=8'd87;
		data_a[16612]<=8'd97;
		data_a[16613]<=8'd110;
		data_a[16614]<=8'd121;
		data_a[16615]<=8'd127;
		data_a[16616]<=8'd128;
		data_a[16617]<=8'd136;
		data_a[16618]<=8'd128;
		data_a[16619]<=8'd123;
		data_a[16620]<=8'd106;
		data_a[16621]<=8'd91;
		data_a[16622]<=8'd91;
		data_a[16623]<=8'd70;
		data_a[16624]<=8'd69;
		data_a[16625]<=8'd57;
		data_a[16626]<=8'd62;
		data_a[16627]<=8'd60;
		data_a[16628]<=8'd64;
		data_a[16629]<=8'd74;
		data_a[16630]<=8'd71;
		data_a[16631]<=8'd95;
		data_a[16632]<=8'd64;
		data_a[16633]<=8'd135;
		data_a[16634]<=8'd235;
		data_a[16635]<=8'd249;
		data_a[16636]<=8'd245;
		data_a[16637]<=8'd245;
		data_a[16638]<=8'd246;
		data_a[16639]<=8'd245;
		data_a[16640]<=8'd247;
		data_a[16641]<=8'd248;
		data_a[16642]<=8'd245;
		data_a[16643]<=8'd247;
		data_a[16644]<=8'd245;
		data_a[16645]<=8'd248;
		data_a[16646]<=8'd248;
		data_a[16647]<=8'd247;
		data_a[16648]<=8'd248;
		data_a[16649]<=8'd247;
		data_a[16650]<=8'd255;
		data_a[16651]<=8'd83;
		data_a[16652]<=8'd83;
		data_a[16653]<=8'd80;
		data_a[16654]<=8'd77;
		data_a[16655]<=8'd76;
		data_a[16656]<=8'd69;
		data_a[16657]<=8'd52;
		data_a[16658]<=8'd55;
		data_a[16659]<=8'd55;
		data_a[16660]<=8'd75;
		data_a[16661]<=8'd73;
		data_a[16662]<=8'd73;
		data_a[16663]<=8'd66;
		data_a[16664]<=8'd72;
		data_a[16665]<=8'd76;
		data_a[16666]<=8'd71;
		data_a[16667]<=8'd69;
		data_a[16668]<=8'd56;
		data_a[16669]<=8'd110;
		data_a[16670]<=8'd58;
		data_a[16671]<=8'd149;
		data_a[16672]<=8'd154;
		data_a[16673]<=8'd157;
		data_a[16674]<=8'd158;
		data_a[16675]<=8'd162;
		data_a[16676]<=8'd164;
		data_a[16677]<=8'd165;
		data_a[16678]<=8'd130;
		data_a[16679]<=8'd108;
		data_a[16680]<=8'd113;
		data_a[16681]<=8'd115;
		data_a[16682]<=8'd113;
		data_a[16683]<=8'd113;
		data_a[16684]<=8'd106;
		data_a[16685]<=8'd85;
		data_a[16686]<=8'd90;
		data_a[16687]<=8'd83;
		data_a[16688]<=8'd89;
		data_a[16689]<=8'd82;
		data_a[16690]<=8'd90;
		data_a[16691]<=8'd94;
		data_a[16692]<=8'd98;
		data_a[16693]<=8'd103;
		data_a[16694]<=8'd100;
		data_a[16695]<=8'd94;
		data_a[16696]<=8'd91;
		data_a[16697]<=8'd79;
		data_a[16698]<=8'd85;
		data_a[16699]<=8'd84;
		data_a[16700]<=8'd86;
		data_a[16701]<=8'd96;
		data_a[16702]<=8'd99;
		data_a[16703]<=8'd96;
		data_a[16704]<=8'd82;
		data_a[16705]<=8'd72;
		data_a[16706]<=8'd76;
		data_a[16707]<=8'd90;
		data_a[16708]<=8'd99;
		data_a[16709]<=8'd111;
		data_a[16710]<=8'd124;
		data_a[16711]<=8'd129;
		data_a[16712]<=8'd141;
		data_a[16713]<=8'd164;
		data_a[16714]<=8'd229;
		data_a[16715]<=8'd230;
		data_a[16716]<=8'd224;
		data_a[16717]<=8'd227;
		data_a[16718]<=8'd233;
		data_a[16719]<=8'd228;
		data_a[16720]<=8'd228;
		data_a[16721]<=8'd234;
		data_a[16722]<=8'd231;
		data_a[16723]<=8'd230;
		data_a[16724]<=8'd234;
		data_a[16725]<=8'd233;
		data_a[16726]<=8'd241;
		data_a[16727]<=8'd242;
		data_a[16728]<=8'd245;
		data_a[16729]<=8'd241;
		data_a[16730]<=8'd242;
		data_a[16731]<=8'd240;
		data_a[16732]<=8'd244;
		data_a[16733]<=8'd237;
		data_a[16734]<=8'd242;
		data_a[16735]<=8'd220;
		data_a[16736]<=8'd80;
		data_a[16737]<=8'd71;
		data_a[16738]<=8'd71;
		data_a[16739]<=8'd71;
		data_a[16740]<=8'd83;
		data_a[16741]<=8'd99;
		data_a[16742]<=8'd120;
		data_a[16743]<=8'd123;
		data_a[16744]<=8'd110;
		data_a[16745]<=8'd86;
		data_a[16746]<=8'd88;
		data_a[16747]<=8'd113;
		data_a[16748]<=8'd118;
		data_a[16749]<=8'd119;
		data_a[16750]<=8'd115;
		data_a[16751]<=8'd119;
		data_a[16752]<=8'd102;
		data_a[16753]<=8'd93;
		data_a[16754]<=8'd87;
		data_a[16755]<=8'd69;
		data_a[16756]<=8'd68;
		data_a[16757]<=8'd67;
		data_a[16758]<=8'd65;
		data_a[16759]<=8'd73;
		data_a[16760]<=8'd71;
		data_a[16761]<=8'd93;
		data_a[16762]<=8'd96;
		data_a[16763]<=8'd105;
		data_a[16764]<=8'd121;
		data_a[16765]<=8'd121;
		data_a[16766]<=8'd132;
		data_a[16767]<=8'd135;
		data_a[16768]<=8'd133;
		data_a[16769]<=8'd123;
		data_a[16770]<=8'd99;
		data_a[16771]<=8'd90;
		data_a[16772]<=8'd79;
		data_a[16773]<=8'd69;
		data_a[16774]<=8'd64;
		data_a[16775]<=8'd58;
		data_a[16776]<=8'd63;
		data_a[16777]<=8'd60;
		data_a[16778]<=8'd58;
		data_a[16779]<=8'd69;
		data_a[16780]<=8'd73;
		data_a[16781]<=8'd75;
		data_a[16782]<=8'd73;
		data_a[16783]<=8'd209;
		data_a[16784]<=8'd253;
		data_a[16785]<=8'd245;
		data_a[16786]<=8'd245;
		data_a[16787]<=8'd245;
		data_a[16788]<=8'd246;
		data_a[16789]<=8'd245;
		data_a[16790]<=8'd248;
		data_a[16791]<=8'd249;
		data_a[16792]<=8'd245;
		data_a[16793]<=8'd247;
		data_a[16794]<=8'd244;
		data_a[16795]<=8'd247;
		data_a[16796]<=8'd246;
		data_a[16797]<=8'd245;
		data_a[16798]<=8'd247;
		data_a[16799]<=8'd247;
		data_a[16800]<=8'd253;
		data_a[16801]<=8'd89;
		data_a[16802]<=8'd84;
		data_a[16803]<=8'd82;
		data_a[16804]<=8'd82;
		data_a[16805]<=8'd83;
		data_a[16806]<=8'd71;
		data_a[16807]<=8'd50;
		data_a[16808]<=8'd58;
		data_a[16809]<=8'd63;
		data_a[16810]<=8'd73;
		data_a[16811]<=8'd72;
		data_a[16812]<=8'd73;
		data_a[16813]<=8'd77;
		data_a[16814]<=8'd83;
		data_a[16815]<=8'd77;
		data_a[16816]<=8'd72;
		data_a[16817]<=8'd69;
		data_a[16818]<=8'd50;
		data_a[16819]<=8'd92;
		data_a[16820]<=8'd50;
		data_a[16821]<=8'd153;
		data_a[16822]<=8'd157;
		data_a[16823]<=8'd157;
		data_a[16824]<=8'd163;
		data_a[16825]<=8'd162;
		data_a[16826]<=8'd165;
		data_a[16827]<=8'd166;
		data_a[16828]<=8'd135;
		data_a[16829]<=8'd113;
		data_a[16830]<=8'd112;
		data_a[16831]<=8'd110;
		data_a[16832]<=8'd108;
		data_a[16833]<=8'd115;
		data_a[16834]<=8'd111;
		data_a[16835]<=8'd88;
		data_a[16836]<=8'd97;
		data_a[16837]<=8'd92;
		data_a[16838]<=8'd56;
		data_a[16839]<=8'd60;
		data_a[16840]<=8'd74;
		data_a[16841]<=8'd84;
		data_a[16842]<=8'd81;
		data_a[16843]<=8'd96;
		data_a[16844]<=8'd93;
		data_a[16845]<=8'd91;
		data_a[16846]<=8'd90;
		data_a[16847]<=8'd79;
		data_a[16848]<=8'd81;
		data_a[16849]<=8'd85;
		data_a[16850]<=8'd82;
		data_a[16851]<=8'd92;
		data_a[16852]<=8'd93;
		data_a[16853]<=8'd107;
		data_a[16854]<=8'd93;
		data_a[16855]<=8'd79;
		data_a[16856]<=8'd74;
		data_a[16857]<=8'd93;
		data_a[16858]<=8'd98;
		data_a[16859]<=8'd116;
		data_a[16860]<=8'd123;
		data_a[16861]<=8'd128;
		data_a[16862]<=8'd131;
		data_a[16863]<=8'd204;
		data_a[16864]<=8'd225;
		data_a[16865]<=8'd224;
		data_a[16866]<=8'd226;
		data_a[16867]<=8'd230;
		data_a[16868]<=8'd231;
		data_a[16869]<=8'd230;
		data_a[16870]<=8'd231;
		data_a[16871]<=8'd234;
		data_a[16872]<=8'd233;
		data_a[16873]<=8'd236;
		data_a[16874]<=8'd230;
		data_a[16875]<=8'd236;
		data_a[16876]<=8'd239;
		data_a[16877]<=8'd246;
		data_a[16878]<=8'd243;
		data_a[16879]<=8'd238;
		data_a[16880]<=8'd237;
		data_a[16881]<=8'd244;
		data_a[16882]<=8'd240;
		data_a[16883]<=8'd240;
		data_a[16884]<=8'd232;
		data_a[16885]<=8'd238;
		data_a[16886]<=8'd149;
		data_a[16887]<=8'd62;
		data_a[16888]<=8'd70;
		data_a[16889]<=8'd69;
		data_a[16890]<=8'd80;
		data_a[16891]<=8'd99;
		data_a[16892]<=8'd114;
		data_a[16893]<=8'd122;
		data_a[16894]<=8'd111;
		data_a[16895]<=8'd94;
		data_a[16896]<=8'd97;
		data_a[16897]<=8'd110;
		data_a[16898]<=8'd121;
		data_a[16899]<=8'd122;
		data_a[16900]<=8'd116;
		data_a[16901]<=8'd107;
		data_a[16902]<=8'd94;
		data_a[16903]<=8'd83;
		data_a[16904]<=8'd77;
		data_a[16905]<=8'd66;
		data_a[16906]<=8'd66;
		data_a[16907]<=8'd70;
		data_a[16908]<=8'd68;
		data_a[16909]<=8'd74;
		data_a[16910]<=8'd74;
		data_a[16911]<=8'd98;
		data_a[16912]<=8'd94;
		data_a[16913]<=8'd105;
		data_a[16914]<=8'd113;
		data_a[16915]<=8'd124;
		data_a[16916]<=8'd141;
		data_a[16917]<=8'd142;
		data_a[16918]<=8'd130;
		data_a[16919]<=8'd119;
		data_a[16920]<=8'd97;
		data_a[16921]<=8'd87;
		data_a[16922]<=8'd74;
		data_a[16923]<=8'd67;
		data_a[16924]<=8'd65;
		data_a[16925]<=8'd56;
		data_a[16926]<=8'd59;
		data_a[16927]<=8'd54;
		data_a[16928]<=8'd54;
		data_a[16929]<=8'd67;
		data_a[16930]<=8'd74;
		data_a[16931]<=8'd96;
		data_a[16932]<=8'd122;
		data_a[16933]<=8'd246;
		data_a[16934]<=8'd243;
		data_a[16935]<=8'd243;
		data_a[16936]<=8'd249;
		data_a[16937]<=8'd246;
		data_a[16938]<=8'd249;
		data_a[16939]<=8'd248;
		data_a[16940]<=8'd248;
		data_a[16941]<=8'd250;
		data_a[16942]<=8'd243;
		data_a[16943]<=8'd247;
		data_a[16944]<=8'd247;
		data_a[16945]<=8'd247;
		data_a[16946]<=8'd247;
		data_a[16947]<=8'd246;
		data_a[16948]<=8'd246;
		data_a[16949]<=8'd246;
		data_a[16950]<=8'd255;
		data_a[16951]<=8'd92;
		data_a[16952]<=8'd88;
		data_a[16953]<=8'd86;
		data_a[16954]<=8'd84;
		data_a[16955]<=8'd83;
		data_a[16956]<=8'd72;
		data_a[16957]<=8'd53;
		data_a[16958]<=8'd58;
		data_a[16959]<=8'd55;
		data_a[16960]<=8'd65;
		data_a[16961]<=8'd74;
		data_a[16962]<=8'd78;
		data_a[16963]<=8'd74;
		data_a[16964]<=8'd73;
		data_a[16965]<=8'd67;
		data_a[16966]<=8'd72;
		data_a[16967]<=8'd69;
		data_a[16968]<=8'd55;
		data_a[16969]<=8'd89;
		data_a[16970]<=8'd50;
		data_a[16971]<=8'd159;
		data_a[16972]<=8'd153;
		data_a[16973]<=8'd156;
		data_a[16974]<=8'd161;
		data_a[16975]<=8'd165;
		data_a[16976]<=8'd164;
		data_a[16977]<=8'd170;
		data_a[16978]<=8'd166;
		data_a[16979]<=8'd116;
		data_a[16980]<=8'd92;
		data_a[16981]<=8'd110;
		data_a[16982]<=8'd116;
		data_a[16983]<=8'd114;
		data_a[16984]<=8'd114;
		data_a[16985]<=8'd93;
		data_a[16986]<=8'd89;
		data_a[16987]<=8'd100;
		data_a[16988]<=8'd85;
		data_a[16989]<=8'd75;
		data_a[16990]<=8'd78;
		data_a[16991]<=8'd90;
		data_a[16992]<=8'd95;
		data_a[16993]<=8'd89;
		data_a[16994]<=8'd82;
		data_a[16995]<=8'd84;
		data_a[16996]<=8'd78;
		data_a[16997]<=8'd88;
		data_a[16998]<=8'd84;
		data_a[16999]<=8'd85;
		data_a[17000]<=8'd83;
		data_a[17001]<=8'd88;
		data_a[17002]<=8'd89;
		data_a[17003]<=8'd80;
		data_a[17004]<=8'd90;
		data_a[17005]<=8'd79;
		data_a[17006]<=8'd79;
		data_a[17007]<=8'd90;
		data_a[17008]<=8'd105;
		data_a[17009]<=8'd118;
		data_a[17010]<=8'd112;
		data_a[17011]<=8'd129;
		data_a[17012]<=8'd154;
		data_a[17013]<=8'd224;
		data_a[17014]<=8'd228;
		data_a[17015]<=8'd228;
		data_a[17016]<=8'd229;
		data_a[17017]<=8'd232;
		data_a[17018]<=8'd232;
		data_a[17019]<=8'd232;
		data_a[17020]<=8'd232;
		data_a[17021]<=8'd234;
		data_a[17022]<=8'd235;
		data_a[17023]<=8'd232;
		data_a[17024]<=8'd236;
		data_a[17025]<=8'd234;
		data_a[17026]<=8'd249;
		data_a[17027]<=8'd245;
		data_a[17028]<=8'd243;
		data_a[17029]<=8'd238;
		data_a[17030]<=8'd241;
		data_a[17031]<=8'd242;
		data_a[17032]<=8'd239;
		data_a[17033]<=8'd240;
		data_a[17034]<=8'd241;
		data_a[17035]<=8'd234;
		data_a[17036]<=8'd215;
		data_a[17037]<=8'd73;
		data_a[17038]<=8'd70;
		data_a[17039]<=8'd69;
		data_a[17040]<=8'd70;
		data_a[17041]<=8'd77;
		data_a[17042]<=8'd100;
		data_a[17043]<=8'd113;
		data_a[17044]<=8'd109;
		data_a[17045]<=8'd103;
		data_a[17046]<=8'd106;
		data_a[17047]<=8'd114;
		data_a[17048]<=8'd120;
		data_a[17049]<=8'd120;
		data_a[17050]<=8'd116;
		data_a[17051]<=8'd109;
		data_a[17052]<=8'd98;
		data_a[17053]<=8'd88;
		data_a[17054]<=8'd76;
		data_a[17055]<=8'd71;
		data_a[17056]<=8'd70;
		data_a[17057]<=8'd70;
		data_a[17058]<=8'd68;
		data_a[17059]<=8'd78;
		data_a[17060]<=8'd77;
		data_a[17061]<=8'd92;
		data_a[17062]<=8'd113;
		data_a[17063]<=8'd115;
		data_a[17064]<=8'd130;
		data_a[17065]<=8'd141;
		data_a[17066]<=8'd134;
		data_a[17067]<=8'd140;
		data_a[17068]<=8'd128;
		data_a[17069]<=8'd108;
		data_a[17070]<=8'd88;
		data_a[17071]<=8'd80;
		data_a[17072]<=8'd71;
		data_a[17073]<=8'd64;
		data_a[17074]<=8'd65;
		data_a[17075]<=8'd48;
		data_a[17076]<=8'd63;
		data_a[17077]<=8'd54;
		data_a[17078]<=8'd54;
		data_a[17079]<=8'd78;
		data_a[17080]<=8'd62;
		data_a[17081]<=8'd106;
		data_a[17082]<=8'd108;
		data_a[17083]<=8'd125;
		data_a[17084]<=8'd140;
		data_a[17085]<=8'd170;
		data_a[17086]<=8'd244;
		data_a[17087]<=8'd252;
		data_a[17088]<=8'd242;
		data_a[17089]<=8'd245;
		data_a[17090]<=8'd242;
		data_a[17091]<=8'd249;
		data_a[17092]<=8'd248;
		data_a[17093]<=8'd243;
		data_a[17094]<=8'd246;
		data_a[17095]<=8'd246;
		data_a[17096]<=8'd246;
		data_a[17097]<=8'd246;
		data_a[17098]<=8'd246;
		data_a[17099]<=8'd245;
		data_a[17100]<=8'd255;
		data_a[17101]<=8'd93;
		data_a[17102]<=8'd91;
		data_a[17103]<=8'd90;
		data_a[17104]<=8'd84;
		data_a[17105]<=8'd81;
		data_a[17106]<=8'd72;
		data_a[17107]<=8'd57;
		data_a[17108]<=8'd55;
		data_a[17109]<=8'd56;
		data_a[17110]<=8'd70;
		data_a[17111]<=8'd78;
		data_a[17112]<=8'd77;
		data_a[17113]<=8'd69;
		data_a[17114]<=8'd73;
		data_a[17115]<=8'd74;
		data_a[17116]<=8'd73;
		data_a[17117]<=8'd71;
		data_a[17118]<=8'd54;
		data_a[17119]<=8'd82;
		data_a[17120]<=8'd39;
		data_a[17121]<=8'd155;
		data_a[17122]<=8'd153;
		data_a[17123]<=8'd160;
		data_a[17124]<=8'd158;
		data_a[17125]<=8'd170;
		data_a[17126]<=8'd168;
		data_a[17127]<=8'd175;
		data_a[17128]<=8'd169;
		data_a[17129]<=8'd102;
		data_a[17130]<=8'd109;
		data_a[17131]<=8'd104;
		data_a[17132]<=8'd117;
		data_a[17133]<=8'd112;
		data_a[17134]<=8'd114;
		data_a[17135]<=8'd100;
		data_a[17136]<=8'd92;
		data_a[17137]<=8'd111;
		data_a[17138]<=8'd113;
		data_a[17139]<=8'd100;
		data_a[17140]<=8'd75;
		data_a[17141]<=8'd89;
		data_a[17142]<=8'd99;
		data_a[17143]<=8'd90;
		data_a[17144]<=8'd96;
		data_a[17145]<=8'd90;
		data_a[17146]<=8'd82;
		data_a[17147]<=8'd88;
		data_a[17148]<=8'd82;
		data_a[17149]<=8'd75;
		data_a[17150]<=8'd78;
		data_a[17151]<=8'd79;
		data_a[17152]<=8'd66;
		data_a[17153]<=8'd61;
		data_a[17154]<=8'd69;
		data_a[17155]<=8'd79;
		data_a[17156]<=8'd87;
		data_a[17157]<=8'd91;
		data_a[17158]<=8'd106;
		data_a[17159]<=8'd117;
		data_a[17160]<=8'd116;
		data_a[17161]<=8'd126;
		data_a[17162]<=8'd195;
		data_a[17163]<=8'd231;
		data_a[17164]<=8'd229;
		data_a[17165]<=8'd230;
		data_a[17166]<=8'd231;
		data_a[17167]<=8'd232;
		data_a[17168]<=8'd233;
		data_a[17169]<=8'd233;
		data_a[17170]<=8'd234;
		data_a[17171]<=8'd235;
		data_a[17172]<=8'd233;
		data_a[17173]<=8'd235;
		data_a[17174]<=8'd231;
		data_a[17175]<=8'd237;
		data_a[17176]<=8'd212;
		data_a[17177]<=8'd244;
		data_a[17178]<=8'd244;
		data_a[17179]<=8'd243;
		data_a[17180]<=8'd240;
		data_a[17181]<=8'd247;
		data_a[17182]<=8'd240;
		data_a[17183]<=8'd238;
		data_a[17184]<=8'd243;
		data_a[17185]<=8'd234;
		data_a[17186]<=8'd235;
		data_a[17187]<=8'd84;
		data_a[17188]<=8'd66;
		data_a[17189]<=8'd68;
		data_a[17190]<=8'd70;
		data_a[17191]<=8'd73;
		data_a[17192]<=8'd94;
		data_a[17193]<=8'd96;
		data_a[17194]<=8'd98;
		data_a[17195]<=8'd115;
		data_a[17196]<=8'd108;
		data_a[17197]<=8'd114;
		data_a[17198]<=8'd119;
		data_a[17199]<=8'd120;
		data_a[17200]<=8'd118;
		data_a[17201]<=8'd111;
		data_a[17202]<=8'd98;
		data_a[17203]<=8'd85;
		data_a[17204]<=8'd78;
		data_a[17205]<=8'd79;
		data_a[17206]<=8'd83;
		data_a[17207]<=8'd79;
		data_a[17208]<=8'd71;
		data_a[17209]<=8'd80;
		data_a[17210]<=8'd91;
		data_a[17211]<=8'd111;
		data_a[17212]<=8'd122;
		data_a[17213]<=8'd125;
		data_a[17214]<=8'd140;
		data_a[17215]<=8'd135;
		data_a[17216]<=8'd138;
		data_a[17217]<=8'd129;
		data_a[17218]<=8'd112;
		data_a[17219]<=8'd93;
		data_a[17220]<=8'd81;
		data_a[17221]<=8'd73;
		data_a[17222]<=8'd77;
		data_a[17223]<=8'd72;
		data_a[17224]<=8'd67;
		data_a[17225]<=8'd61;
		data_a[17226]<=8'd55;
		data_a[17227]<=8'd56;
		data_a[17228]<=8'd65;
		data_a[17229]<=8'd59;
		data_a[17230]<=8'd68;
		data_a[17231]<=8'd104;
		data_a[17232]<=8'd155;
		data_a[17233]<=8'd100;
		data_a[17234]<=8'd114;
		data_a[17235]<=8'd125;
		data_a[17236]<=8'd132;
		data_a[17237]<=8'd242;
		data_a[17238]<=8'd243;
		data_a[17239]<=8'd246;
		data_a[17240]<=8'd246;
		data_a[17241]<=8'd241;
		data_a[17242]<=8'd249;
		data_a[17243]<=8'd245;
		data_a[17244]<=8'd245;
		data_a[17245]<=8'd245;
		data_a[17246]<=8'd245;
		data_a[17247]<=8'd245;
		data_a[17248]<=8'd245;
		data_a[17249]<=8'd244;
		data_a[17250]<=8'd254;
		data_a[17251]<=8'd92;
		data_a[17252]<=8'd91;
		data_a[17253]<=8'd91;
		data_a[17254]<=8'd86;
		data_a[17255]<=8'd81;
		data_a[17256]<=8'd73;
		data_a[17257]<=8'd61;
		data_a[17258]<=8'd52;
		data_a[17259]<=8'd55;
		data_a[17260]<=8'd68;
		data_a[17261]<=8'd72;
		data_a[17262]<=8'd74;
		data_a[17263]<=8'd74;
		data_a[17264]<=8'd77;
		data_a[17265]<=8'd71;
		data_a[17266]<=8'd73;
		data_a[17267]<=8'd72;
		data_a[17268]<=8'd52;
		data_a[17269]<=8'd120;
		data_a[17270]<=8'd49;
		data_a[17271]<=8'd155;
		data_a[17272]<=8'd161;
		data_a[17273]<=8'd159;
		data_a[17274]<=8'd164;
		data_a[17275]<=8'd161;
		data_a[17276]<=8'd168;
		data_a[17277]<=8'd173;
		data_a[17278]<=8'd175;
		data_a[17279]<=8'd119;
		data_a[17280]<=8'd106;
		data_a[17281]<=8'd103;
		data_a[17282]<=8'd116;
		data_a[17283]<=8'd115;
		data_a[17284]<=8'd111;
		data_a[17285]<=8'd104;
		data_a[17286]<=8'd99;
		data_a[17287]<=8'd106;
		data_a[17288]<=8'd108;
		data_a[17289]<=8'd107;
		data_a[17290]<=8'd105;
		data_a[17291]<=8'd86;
		data_a[17292]<=8'd102;
		data_a[17293]<=8'd111;
		data_a[17294]<=8'd101;
		data_a[17295]<=8'd104;
		data_a[17296]<=8'd82;
		data_a[17297]<=8'd96;
		data_a[17298]<=8'd85;
		data_a[17299]<=8'd88;
		data_a[17300]<=8'd89;
		data_a[17301]<=8'd90;
		data_a[17302]<=8'd60;
		data_a[17303]<=8'd56;
		data_a[17304]<=8'd68;
		data_a[17305]<=8'd87;
		data_a[17306]<=8'd89;
		data_a[17307]<=8'd93;
		data_a[17308]<=8'd109;
		data_a[17309]<=8'd123;
		data_a[17310]<=8'd111;
		data_a[17311]<=8'd138;
		data_a[17312]<=8'd211;
		data_a[17313]<=8'd233;
		data_a[17314]<=8'd228;
		data_a[17315]<=8'd230;
		data_a[17316]<=8'd232;
		data_a[17317]<=8'd232;
		data_a[17318]<=8'd233;
		data_a[17319]<=8'd235;
		data_a[17320]<=8'd236;
		data_a[17321]<=8'd235;
		data_a[17322]<=8'd237;
		data_a[17323]<=8'd233;
		data_a[17324]<=8'd234;
		data_a[17325]<=8'd235;
		data_a[17326]<=8'd214;
		data_a[17327]<=8'd248;
		data_a[17328]<=8'd248;
		data_a[17329]<=8'd239;
		data_a[17330]<=8'd244;
		data_a[17331]<=8'd241;
		data_a[17332]<=8'd239;
		data_a[17333]<=8'd240;
		data_a[17334]<=8'd248;
		data_a[17335]<=8'd239;
		data_a[17336]<=8'd249;
		data_a[17337]<=8'd75;
		data_a[17338]<=8'd73;
		data_a[17339]<=8'd68;
		data_a[17340]<=8'd64;
		data_a[17341]<=8'd66;
		data_a[17342]<=8'd84;
		data_a[17343]<=8'd92;
		data_a[17344]<=8'd95;
		data_a[17345]<=8'd113;
		data_a[17346]<=8'd107;
		data_a[17347]<=8'd112;
		data_a[17348]<=8'd117;
		data_a[17349]<=8'd120;
		data_a[17350]<=8'd120;
		data_a[17351]<=8'd114;
		data_a[17352]<=8'd101;
		data_a[17353]<=8'd89;
		data_a[17354]<=8'd85;
		data_a[17355]<=8'd74;
		data_a[17356]<=8'd84;
		data_a[17357]<=8'd77;
		data_a[17358]<=8'd89;
		data_a[17359]<=8'd82;
		data_a[17360]<=8'd106;
		data_a[17361]<=8'd121;
		data_a[17362]<=8'd133;
		data_a[17363]<=8'd137;
		data_a[17364]<=8'd136;
		data_a[17365]<=8'd144;
		data_a[17366]<=8'd133;
		data_a[17367]<=8'd128;
		data_a[17368]<=8'd105;
		data_a[17369]<=8'd86;
		data_a[17370]<=8'd79;
		data_a[17371]<=8'd68;
		data_a[17372]<=8'd68;
		data_a[17373]<=8'd60;
		data_a[17374]<=8'd60;
		data_a[17375]<=8'd59;
		data_a[17376]<=8'd48;
		data_a[17377]<=8'd57;
		data_a[17378]<=8'd55;
		data_a[17379]<=8'd62;
		data_a[17380]<=8'd67;
		data_a[17381]<=8'd113;
		data_a[17382]<=8'd181;
		data_a[17383]<=8'd70;
		data_a[17384]<=8'd85;
		data_a[17385]<=8'd103;
		data_a[17386]<=8'd127;
		data_a[17387]<=8'd150;
		data_a[17388]<=8'd248;
		data_a[17389]<=8'd244;
		data_a[17390]<=8'd248;
		data_a[17391]<=8'd247;
		data_a[17392]<=8'd240;
		data_a[17393]<=8'd244;
		data_a[17394]<=8'd244;
		data_a[17395]<=8'd244;
		data_a[17396]<=8'd244;
		data_a[17397]<=8'd244;
		data_a[17398]<=8'd244;
		data_a[17399]<=8'd244;
		data_a[17400]<=8'd255;
		data_a[17401]<=8'd92;
		data_a[17402]<=8'd91;
		data_a[17403]<=8'd92;
		data_a[17404]<=8'd87;
		data_a[17405]<=8'd82;
		data_a[17406]<=8'd74;
		data_a[17407]<=8'd62;
		data_a[17408]<=8'd46;
		data_a[17409]<=8'd58;
		data_a[17410]<=8'd75;
		data_a[17411]<=8'd76;
		data_a[17412]<=8'd72;
		data_a[17413]<=8'd71;
		data_a[17414]<=8'd76;
		data_a[17415]<=8'd72;
		data_a[17416]<=8'd70;
		data_a[17417]<=8'd70;
		data_a[17418]<=8'd71;
		data_a[17419]<=8'd71;
		data_a[17420]<=8'd47;
		data_a[17421]<=8'd160;
		data_a[17422]<=8'd155;
		data_a[17423]<=8'd164;
		data_a[17424]<=8'd163;
		data_a[17425]<=8'd172;
		data_a[17426]<=8'd170;
		data_a[17427]<=8'd177;
		data_a[17428]<=8'd158;
		data_a[17429]<=8'd152;
		data_a[17430]<=8'd107;
		data_a[17431]<=8'd99;
		data_a[17432]<=8'd114;
		data_a[17433]<=8'd116;
		data_a[17434]<=8'd111;
		data_a[17435]<=8'd109;
		data_a[17436]<=8'd103;
		data_a[17437]<=8'd107;
		data_a[17438]<=8'd108;
		data_a[17439]<=8'd113;
		data_a[17440]<=8'd103;
		data_a[17441]<=8'd122;
		data_a[17442]<=8'd88;
		data_a[17443]<=8'd100;
		data_a[17444]<=8'd97;
		data_a[17445]<=8'd121;
		data_a[17446]<=8'd94;
		data_a[17447]<=8'd110;
		data_a[17448]<=8'd100;
		data_a[17449]<=8'd105;
		data_a[17450]<=8'd78;
		data_a[17451]<=8'd82;
		data_a[17452]<=8'd69;
		data_a[17453]<=8'd64;
		data_a[17454]<=8'd94;
		data_a[17455]<=8'd89;
		data_a[17456]<=8'd80;
		data_a[17457]<=8'd104;
		data_a[17458]<=8'd114;
		data_a[17459]<=8'd120;
		data_a[17460]<=8'd117;
		data_a[17461]<=8'd127;
		data_a[17462]<=8'd229;
		data_a[17463]<=8'd230;
		data_a[17464]<=8'd230;
		data_a[17465]<=8'd232;
		data_a[17466]<=8'd233;
		data_a[17467]<=8'd233;
		data_a[17468]<=8'd234;
		data_a[17469]<=8'd235;
		data_a[17470]<=8'd236;
		data_a[17471]<=8'd236;
		data_a[17472]<=8'd238;
		data_a[17473]<=8'd233;
		data_a[17474]<=8'd237;
		data_a[17475]<=8'd233;
		data_a[17476]<=8'd238;
		data_a[17477]<=8'd246;
		data_a[17478]<=8'd241;
		data_a[17479]<=8'd244;
		data_a[17480]<=8'd243;
		data_a[17481]<=8'd238;
		data_a[17482]<=8'd243;
		data_a[17483]<=8'd243;
		data_a[17484]<=8'd237;
		data_a[17485]<=8'd245;
		data_a[17486]<=8'd199;
		data_a[17487]<=8'd50;
		data_a[17488]<=8'd67;
		data_a[17489]<=8'd68;
		data_a[17490]<=8'd72;
		data_a[17491]<=8'd66;
		data_a[17492]<=8'd65;
		data_a[17493]<=8'd83;
		data_a[17494]<=8'd93;
		data_a[17495]<=8'd104;
		data_a[17496]<=8'd107;
		data_a[17497]<=8'd111;
		data_a[17498]<=8'd114;
		data_a[17499]<=8'd117;
		data_a[17500]<=8'd118;
		data_a[17501]<=8'd117;
		data_a[17502]<=8'd112;
		data_a[17503]<=8'd106;
		data_a[17504]<=8'd95;
		data_a[17505]<=8'd93;
		data_a[17506]<=8'd86;
		data_a[17507]<=8'd107;
		data_a[17508]<=8'd97;
		data_a[17509]<=8'd108;
		data_a[17510]<=8'd112;
		data_a[17511]<=8'd128;
		data_a[17512]<=8'd129;
		data_a[17513]<=8'd136;
		data_a[17514]<=8'd126;
		data_a[17515]<=8'd120;
		data_a[17516]<=8'd127;
		data_a[17517]<=8'd103;
		data_a[17518]<=8'd91;
		data_a[17519]<=8'd78;
		data_a[17520]<=8'd70;
		data_a[17521]<=8'd69;
		data_a[17522]<=8'd61;
		data_a[17523]<=8'd57;
		data_a[17524]<=8'd76;
		data_a[17525]<=8'd53;
		data_a[17526]<=8'd57;
		data_a[17527]<=8'd50;
		data_a[17528]<=8'd59;
		data_a[17529]<=8'd58;
		data_a[17530]<=8'd72;
		data_a[17531]<=8'd115;
		data_a[17532]<=8'd160;
		data_a[17533]<=8'd69;
		data_a[17534]<=8'd81;
		data_a[17535]<=8'd94;
		data_a[17536]<=8'd115;
		data_a[17537]<=8'd136;
		data_a[17538]<=8'd164;
		data_a[17539]<=8'd245;
		data_a[17540]<=8'd239;
		data_a[17541]<=8'd248;
		data_a[17542]<=8'd244;
		data_a[17543]<=8'd249;
		data_a[17544]<=8'd244;
		data_a[17545]<=8'd244;
		data_a[17546]<=8'd244;
		data_a[17547]<=8'd244;
		data_a[17548]<=8'd243;
		data_a[17549]<=8'd243;
		data_a[17550]<=8'd255;
		data_a[17551]<=8'd92;
		data_a[17552]<=8'd91;
		data_a[17553]<=8'd91;
		data_a[17554]<=8'd86;
		data_a[17555]<=8'd82;
		data_a[17556]<=8'd73;
		data_a[17557]<=8'd60;
		data_a[17558]<=8'd62;
		data_a[17559]<=8'd61;
		data_a[17560]<=8'd69;
		data_a[17561]<=8'd74;
		data_a[17562]<=8'd79;
		data_a[17563]<=8'd78;
		data_a[17564]<=8'd77;
		data_a[17565]<=8'd69;
		data_a[17566]<=8'd77;
		data_a[17567]<=8'd67;
		data_a[17568]<=8'd54;
		data_a[17569]<=8'd87;
		data_a[17570]<=8'd51;
		data_a[17571]<=8'd158;
		data_a[17572]<=8'd162;
		data_a[17573]<=8'd162;
		data_a[17574]<=8'd171;
		data_a[17575]<=8'd169;
		data_a[17576]<=8'd173;
		data_a[17577]<=8'd179;
		data_a[17578]<=8'd171;
		data_a[17579]<=8'd151;
		data_a[17580]<=8'd102;
		data_a[17581]<=8'd100;
		data_a[17582]<=8'd110;
		data_a[17583]<=8'd111;
		data_a[17584]<=8'd112;
		data_a[17585]<=8'd110;
		data_a[17586]<=8'd99;
		data_a[17587]<=8'd113;
		data_a[17588]<=8'd121;
		data_a[17589]<=8'd120;
		data_a[17590]<=8'd101;
		data_a[17591]<=8'd99;
		data_a[17592]<=8'd102;
		data_a[17593]<=8'd114;
		data_a[17594]<=8'd95;
		data_a[17595]<=8'd98;
		data_a[17596]<=8'd86;
		data_a[17597]<=8'd112;
		data_a[17598]<=8'd93;
		data_a[17599]<=8'd98;
		data_a[17600]<=8'd64;
		data_a[17601]<=8'd78;
		data_a[17602]<=8'd78;
		data_a[17603]<=8'd91;
		data_a[17604]<=8'd104;
		data_a[17605]<=8'd89;
		data_a[17606]<=8'd80;
		data_a[17607]<=8'd106;
		data_a[17608]<=8'd114;
		data_a[17609]<=8'd117;
		data_a[17610]<=8'd107;
		data_a[17611]<=8'd152;
		data_a[17612]<=8'd223;
		data_a[17613]<=8'd234;
		data_a[17614]<=8'd232;
		data_a[17615]<=8'd232;
		data_a[17616]<=8'd233;
		data_a[17617]<=8'd234;
		data_a[17618]<=8'd234;
		data_a[17619]<=8'd234;
		data_a[17620]<=8'd234;
		data_a[17621]<=8'd235;
		data_a[17622]<=8'd235;
		data_a[17623]<=8'd237;
		data_a[17624]<=8'd233;
		data_a[17625]<=8'd235;
		data_a[17626]<=8'd230;
		data_a[17627]<=8'd244;
		data_a[17628]<=8'd239;
		data_a[17629]<=8'd246;
		data_a[17630]<=8'd242;
		data_a[17631]<=8'd236;
		data_a[17632]<=8'd242;
		data_a[17633]<=8'd243;
		data_a[17634]<=8'd245;
		data_a[17635]<=8'd241;
		data_a[17636]<=8'd250;
		data_a[17637]<=8'd171;
		data_a[17638]<=8'd90;
		data_a[17639]<=8'd66;
		data_a[17640]<=8'd67;
		data_a[17641]<=8'd66;
		data_a[17642]<=8'd65;
		data_a[17643]<=8'd83;
		data_a[17644]<=8'd90;
		data_a[17645]<=8'd87;
		data_a[17646]<=8'd103;
		data_a[17647]<=8'd107;
		data_a[17648]<=8'd113;
		data_a[17649]<=8'd117;
		data_a[17650]<=8'd118;
		data_a[17651]<=8'd117;
		data_a[17652]<=8'd115;
		data_a[17653]<=8'd114;
		data_a[17654]<=8'd108;
		data_a[17655]<=8'd107;
		data_a[17656]<=8'd108;
		data_a[17657]<=8'd110;
		data_a[17658]<=8'd109;
		data_a[17659]<=8'd106;
		data_a[17660]<=8'd120;
		data_a[17661]<=8'd121;
		data_a[17662]<=8'd131;
		data_a[17663]<=8'd125;
		data_a[17664]<=8'd116;
		data_a[17665]<=8'd121;
		data_a[17666]<=8'd98;
		data_a[17667]<=8'd93;
		data_a[17668]<=8'd92;
		data_a[17669]<=8'd75;
		data_a[17670]<=8'd73;
		data_a[17671]<=8'd65;
		data_a[17672]<=8'd54;
		data_a[17673]<=8'd51;
		data_a[17674]<=8'd63;
		data_a[17675]<=8'd52;
		data_a[17676]<=8'd55;
		data_a[17677]<=8'd52;
		data_a[17678]<=8'd55;
		data_a[17679]<=8'd60;
		data_a[17680]<=8'd76;
		data_a[17681]<=8'd138;
		data_a[17682]<=8'd172;
		data_a[17683]<=8'd96;
		data_a[17684]<=8'd66;
		data_a[17685]<=8'd87;
		data_a[17686]<=8'd104;
		data_a[17687]<=8'd111;
		data_a[17688]<=8'd148;
		data_a[17689]<=8'd235;
		data_a[17690]<=8'd242;
		data_a[17691]<=8'd243;
		data_a[17692]<=8'd244;
		data_a[17693]<=8'd239;
		data_a[17694]<=8'd244;
		data_a[17695]<=8'd244;
		data_a[17696]<=8'd244;
		data_a[17697]<=8'd244;
		data_a[17698]<=8'd243;
		data_a[17699]<=8'd243;
		data_a[17700]<=8'd254;
		data_a[17701]<=8'd92;
		data_a[17702]<=8'd91;
		data_a[17703]<=8'd90;
		data_a[17704]<=8'd85;
		data_a[17705]<=8'd82;
		data_a[17706]<=8'd74;
		data_a[17707]<=8'd60;
		data_a[17708]<=8'd62;
		data_a[17709]<=8'd61;
		data_a[17710]<=8'd71;
		data_a[17711]<=8'd74;
		data_a[17712]<=8'd73;
		data_a[17713]<=8'd70;
		data_a[17714]<=8'd74;
		data_a[17715]<=8'd73;
		data_a[17716]<=8'd74;
		data_a[17717]<=8'd68;
		data_a[17718]<=8'd57;
		data_a[17719]<=8'd83;
		data_a[17720]<=8'd57;
		data_a[17721]<=8'd162;
		data_a[17722]<=8'd163;
		data_a[17723]<=8'd161;
		data_a[17724]<=8'd163;
		data_a[17725]<=8'd178;
		data_a[17726]<=8'd171;
		data_a[17727]<=8'd179;
		data_a[17728]<=8'd177;
		data_a[17729]<=8'd188;
		data_a[17730]<=8'd77;
		data_a[17731]<=8'd95;
		data_a[17732]<=8'd108;
		data_a[17733]<=8'd107;
		data_a[17734]<=8'd110;
		data_a[17735]<=8'd106;
		data_a[17736]<=8'd92;
		data_a[17737]<=8'd112;
		data_a[17738]<=8'd119;
		data_a[17739]<=8'd113;
		data_a[17740]<=8'd116;
		data_a[17741]<=8'd101;
		data_a[17742]<=8'd103;
		data_a[17743]<=8'd106;
		data_a[17744]<=8'd111;
		data_a[17745]<=8'd94;
		data_a[17746]<=8'd85;
		data_a[17747]<=8'd83;
		data_a[17748]<=8'd83;
		data_a[17749]<=8'd97;
		data_a[17750]<=8'd87;
		data_a[17751]<=8'd101;
		data_a[17752]<=8'd95;
		data_a[17753]<=8'd112;
		data_a[17754]<=8'd100;
		data_a[17755]<=8'd98;
		data_a[17756]<=8'd88;
		data_a[17757]<=8'd106;
		data_a[17758]<=8'd110;
		data_a[17759]<=8'd109;
		data_a[17760]<=8'd116;
		data_a[17761]<=8'd176;
		data_a[17762]<=8'd230;
		data_a[17763]<=8'd230;
		data_a[17764]<=8'd232;
		data_a[17765]<=8'd232;
		data_a[17766]<=8'd233;
		data_a[17767]<=8'd234;
		data_a[17768]<=8'd235;
		data_a[17769]<=8'd233;
		data_a[17770]<=8'd233;
		data_a[17771]<=8'd235;
		data_a[17772]<=8'd236;
		data_a[17773]<=8'd234;
		data_a[17774]<=8'd235;
		data_a[17775]<=8'd236;
		data_a[17776]<=8'd233;
		data_a[17777]<=8'd247;
		data_a[17778]<=8'd248;
		data_a[17779]<=8'd235;
		data_a[17780]<=8'd239;
		data_a[17781]<=8'd245;
		data_a[17782]<=8'd244;
		data_a[17783]<=8'd241;
		data_a[17784]<=8'd243;
		data_a[17785]<=8'd240;
		data_a[17786]<=8'd247;
		data_a[17787]<=8'd253;
		data_a[17788]<=8'd122;
		data_a[17789]<=8'd70;
		data_a[17790]<=8'd66;
		data_a[17791]<=8'd64;
		data_a[17792]<=8'd64;
		data_a[17793]<=8'd69;
		data_a[17794]<=8'd86;
		data_a[17795]<=8'd92;
		data_a[17796]<=8'd95;
		data_a[17797]<=8'd103;
		data_a[17798]<=8'd113;
		data_a[17799]<=8'd120;
		data_a[17800]<=8'd121;
		data_a[17801]<=8'd119;
		data_a[17802]<=8'd116;
		data_a[17803]<=8'd115;
		data_a[17804]<=8'd127;
		data_a[17805]<=8'd123;
		data_a[17806]<=8'd118;
		data_a[17807]<=8'd117;
		data_a[17808]<=8'd119;
		data_a[17809]<=8'd116;
		data_a[17810]<=8'd125;
		data_a[17811]<=8'd111;
		data_a[17812]<=8'd124;
		data_a[17813]<=8'd117;
		data_a[17814]<=8'd113;
		data_a[17815]<=8'd99;
		data_a[17816]<=8'd93;
		data_a[17817]<=8'd88;
		data_a[17818]<=8'd84;
		data_a[17819]<=8'd73;
		data_a[17820]<=8'd72;
		data_a[17821]<=8'd56;
		data_a[17822]<=8'd61;
		data_a[17823]<=8'd66;
		data_a[17824]<=8'd55;
		data_a[17825]<=8'd63;
		data_a[17826]<=8'd50;
		data_a[17827]<=8'd53;
		data_a[17828]<=8'd64;
		data_a[17829]<=8'd61;
		data_a[17830]<=8'd86;
		data_a[17831]<=8'd140;
		data_a[17832]<=8'd150;
		data_a[17833]<=8'd151;
		data_a[17834]<=8'd69;
		data_a[17835]<=8'd82;
		data_a[17836]<=8'd94;
		data_a[17837]<=8'd117;
		data_a[17838]<=8'd127;
		data_a[17839]<=8'd139;
		data_a[17840]<=8'd241;
		data_a[17841]<=8'd244;
		data_a[17842]<=8'd247;
		data_a[17843]<=8'd245;
		data_a[17844]<=8'd244;
		data_a[17845]<=8'd244;
		data_a[17846]<=8'd244;
		data_a[17847]<=8'd244;
		data_a[17848]<=8'd244;
		data_a[17849]<=8'd243;
		data_a[17850]<=8'd254;
		data_a[17851]<=8'd93;
		data_a[17852]<=8'd92;
		data_a[17853]<=8'd91;
		data_a[17854]<=8'd86;
		data_a[17855]<=8'd84;
		data_a[17856]<=8'd76;
		data_a[17857]<=8'd62;
		data_a[17858]<=8'd56;
		data_a[17859]<=8'd60;
		data_a[17860]<=8'd73;
		data_a[17861]<=8'd76;
		data_a[17862]<=8'd75;
		data_a[17863]<=8'd72;
		data_a[17864]<=8'd75;
		data_a[17865]<=8'd72;
		data_a[17866]<=8'd72;
		data_a[17867]<=8'd69;
		data_a[17868]<=8'd61;
		data_a[17869]<=8'd73;
		data_a[17870]<=8'd54;
		data_a[17871]<=8'd162;
		data_a[17872]<=8'd159;
		data_a[17873]<=8'd166;
		data_a[17874]<=8'd167;
		data_a[17875]<=8'd172;
		data_a[17876]<=8'd175;
		data_a[17877]<=8'd180;
		data_a[17878]<=8'd181;
		data_a[17879]<=8'd177;
		data_a[17880]<=8'd91;
		data_a[17881]<=8'd95;
		data_a[17882]<=8'd104;
		data_a[17883]<=8'd106;
		data_a[17884]<=8'd108;
		data_a[17885]<=8'd106;
		data_a[17886]<=8'd97;
		data_a[17887]<=8'd116;
		data_a[17888]<=8'd116;
		data_a[17889]<=8'd115;
		data_a[17890]<=8'd116;
		data_a[17891]<=8'd101;
		data_a[17892]<=8'd103;
		data_a[17893]<=8'd100;
		data_a[17894]<=8'd104;
		data_a[17895]<=8'd105;
		data_a[17896]<=8'd101;
		data_a[17897]<=8'd119;
		data_a[17898]<=8'd106;
		data_a[17899]<=8'd111;
		data_a[17900]<=8'd96;
		data_a[17901]<=8'd98;
		data_a[17902]<=8'd103;
		data_a[17903]<=8'd104;
		data_a[17904]<=8'd102;
		data_a[17905]<=8'd96;
		data_a[17906]<=8'd94;
		data_a[17907]<=8'd102;
		data_a[17908]<=8'd112;
		data_a[17909]<=8'd111;
		data_a[17910]<=8'd116;
		data_a[17911]<=8'd203;
		data_a[17912]<=8'd227;
		data_a[17913]<=8'd231;
		data_a[17914]<=8'd234;
		data_a[17915]<=8'd232;
		data_a[17916]<=8'd233;
		data_a[17917]<=8'd236;
		data_a[17918]<=8'd237;
		data_a[17919]<=8'd235;
		data_a[17920]<=8'd235;
		data_a[17921]<=8'd238;
		data_a[17922]<=8'd233;
		data_a[17923]<=8'd238;
		data_a[17924]<=8'd235;
		data_a[17925]<=8'd239;
		data_a[17926]<=8'd235;
		data_a[17927]<=8'd241;
		data_a[17928]<=8'd243;
		data_a[17929]<=8'd243;
		data_a[17930]<=8'd243;
		data_a[17931]<=8'd241;
		data_a[17932]<=8'd245;
		data_a[17933]<=8'd243;
		data_a[17934]<=8'd242;
		data_a[17935]<=8'd243;
		data_a[17936]<=8'd242;
		data_a[17937]<=8'd239;
		data_a[17938]<=8'd136;
		data_a[17939]<=8'd70;
		data_a[17940]<=8'd64;
		data_a[17941]<=8'd58;
		data_a[17942]<=8'd70;
		data_a[17943]<=8'd71;
		data_a[17944]<=8'd86;
		data_a[17945]<=8'd85;
		data_a[17946]<=8'd91;
		data_a[17947]<=8'd101;
		data_a[17948]<=8'd114;
		data_a[17949]<=8'd123;
		data_a[17950]<=8'd125;
		data_a[17951]<=8'd123;
		data_a[17952]<=8'd122;
		data_a[17953]<=8'd122;
		data_a[17954]<=8'd123;
		data_a[17955]<=8'd124;
		data_a[17956]<=8'd124;
		data_a[17957]<=8'd124;
		data_a[17958]<=8'd121;
		data_a[17959]<=8'd112;
		data_a[17960]<=8'd120;
		data_a[17961]<=8'd105;
		data_a[17962]<=8'd119;
		data_a[17963]<=8'd112;
		data_a[17964]<=8'd107;
		data_a[17965]<=8'd89;
		data_a[17966]<=8'd87;
		data_a[17967]<=8'd93;
		data_a[17968]<=8'd73;
		data_a[17969]<=8'd64;
		data_a[17970]<=8'd65;
		data_a[17971]<=8'd47;
		data_a[17972]<=8'd55;
		data_a[17973]<=8'd64;
		data_a[17974]<=8'd46;
		data_a[17975]<=8'd52;
		data_a[17976]<=8'd55;
		data_a[17977]<=8'd50;
		data_a[17978]<=8'd53;
		data_a[17979]<=8'd69;
		data_a[17980]<=8'd95;
		data_a[17981]<=8'd144;
		data_a[17982]<=8'd157;
		data_a[17983]<=8'd148;
		data_a[17984]<=8'd68;
		data_a[17985]<=8'd74;
		data_a[17986]<=8'd90;
		data_a[17987]<=8'd95;
		data_a[17988]<=8'd119;
		data_a[17989]<=8'd141;
		data_a[17990]<=8'd249;
		data_a[17991]<=8'd246;
		data_a[17992]<=8'd242;
		data_a[17993]<=8'd244;
		data_a[17994]<=8'd244;
		data_a[17995]<=8'd244;
		data_a[17996]<=8'd244;
		data_a[17997]<=8'd244;
		data_a[17998]<=8'd244;
		data_a[17999]<=8'd243;
		data_a[18000]<=8'd253;
		data_a[18001]<=8'd98;
		data_a[18002]<=8'd89;
		data_a[18003]<=8'd91;
		data_a[18004]<=8'd86;
		data_a[18005]<=8'd82;
		data_a[18006]<=8'd71;
		data_a[18007]<=8'd69;
		data_a[18008]<=8'd59;
		data_a[18009]<=8'd64;
		data_a[18010]<=8'd81;
		data_a[18011]<=8'd74;
		data_a[18012]<=8'd77;
		data_a[18013]<=8'd75;
		data_a[18014]<=8'd77;
		data_a[18015]<=8'd70;
		data_a[18016]<=8'd73;
		data_a[18017]<=8'd67;
		data_a[18018]<=8'd67;
		data_a[18019]<=8'd70;
		data_a[18020]<=8'd51;
		data_a[18021]<=8'd162;
		data_a[18022]<=8'd164;
		data_a[18023]<=8'd166;
		data_a[18024]<=8'd166;
		data_a[18025]<=8'd171;
		data_a[18026]<=8'd177;
		data_a[18027]<=8'd180;
		data_a[18028]<=8'd184;
		data_a[18029]<=8'd190;
		data_a[18030]<=8'd123;
		data_a[18031]<=8'd97;
		data_a[18032]<=8'd101;
		data_a[18033]<=8'd102;
		data_a[18034]<=8'd104;
		data_a[18035]<=8'd109;
		data_a[18036]<=8'd102;
		data_a[18037]<=8'd112;
		data_a[18038]<=8'd120;
		data_a[18039]<=8'd116;
		data_a[18040]<=8'd116;
		data_a[18041]<=8'd119;
		data_a[18042]<=8'd96;
		data_a[18043]<=8'd99;
		data_a[18044]<=8'd107;
		data_a[18045]<=8'd104;
		data_a[18046]<=8'd104;
		data_a[18047]<=8'd108;
		data_a[18048]<=8'd110;
		data_a[18049]<=8'd99;
		data_a[18050]<=8'd97;
		data_a[18051]<=8'd101;
		data_a[18052]<=8'd111;
		data_a[18053]<=8'd102;
		data_a[18054]<=8'd97;
		data_a[18055]<=8'd97;
		data_a[18056]<=8'd96;
		data_a[18057]<=8'd99;
		data_a[18058]<=8'd111;
		data_a[18059]<=8'd105;
		data_a[18060]<=8'd133;
		data_a[18061]<=8'd229;
		data_a[18062]<=8'd226;
		data_a[18063]<=8'd233;
		data_a[18064]<=8'd231;
		data_a[18065]<=8'd234;
		data_a[18066]<=8'd236;
		data_a[18067]<=8'd236;
		data_a[18068]<=8'd234;
		data_a[18069]<=8'd233;
		data_a[18070]<=8'd235;
		data_a[18071]<=8'd238;
		data_a[18072]<=8'd235;
		data_a[18073]<=8'd235;
		data_a[18074]<=8'd234;
		data_a[18075]<=8'd233;
		data_a[18076]<=8'd236;
		data_a[18077]<=8'd242;
		data_a[18078]<=8'd244;
		data_a[18079]<=8'd243;
		data_a[18080]<=8'd245;
		data_a[18081]<=8'd244;
		data_a[18082]<=8'd241;
		data_a[18083]<=8'd246;
		data_a[18084]<=8'd244;
		data_a[18085]<=8'd244;
		data_a[18086]<=8'd242;
		data_a[18087]<=8'd244;
		data_a[18088]<=8'd233;
		data_a[18089]<=8'd111;
		data_a[18090]<=8'd57;
		data_a[18091]<=8'd58;
		data_a[18092]<=8'd59;
		data_a[18093]<=8'd67;
		data_a[18094]<=8'd79;
		data_a[18095]<=8'd87;
		data_a[18096]<=8'd85;
		data_a[18097]<=8'd99;
		data_a[18098]<=8'd103;
		data_a[18099]<=8'd117;
		data_a[18100]<=8'd120;
		data_a[18101]<=8'd126;
		data_a[18102]<=8'd129;
		data_a[18103]<=8'd125;
		data_a[18104]<=8'd129;
		data_a[18105]<=8'd117;
		data_a[18106]<=8'd110;
		data_a[18107]<=8'd126;
		data_a[18108]<=8'd116;
		data_a[18109]<=8'd111;
		data_a[18110]<=8'd103;
		data_a[18111]<=8'd99;
		data_a[18112]<=8'd105;
		data_a[18113]<=8'd97;
		data_a[18114]<=8'd91;
		data_a[18115]<=8'd84;
		data_a[18116]<=8'd84;
		data_a[18117]<=8'd74;
		data_a[18118]<=8'd69;
		data_a[18119]<=8'd58;
		data_a[18120]<=8'd50;
		data_a[18121]<=8'd57;
		data_a[18122]<=8'd52;
		data_a[18123]<=8'd53;
		data_a[18124]<=8'd53;
		data_a[18125]<=8'd45;
		data_a[18126]<=8'd52;
		data_a[18127]<=8'd56;
		data_a[18128]<=8'd53;
		data_a[18129]<=8'd72;
		data_a[18130]<=8'd111;
		data_a[18131]<=8'd142;
		data_a[18132]<=8'd157;
		data_a[18133]<=8'd145;
		data_a[18134]<=8'd56;
		data_a[18135]<=8'd70;
		data_a[18136]<=8'd88;
		data_a[18137]<=8'd106;
		data_a[18138]<=8'd120;
		data_a[18139]<=8'd128;
		data_a[18140]<=8'd194;
		data_a[18141]<=8'd250;
		data_a[18142]<=8'd244;
		data_a[18143]<=8'd246;
		data_a[18144]<=8'd242;
		data_a[18145]<=8'd245;
		data_a[18146]<=8'd245;
		data_a[18147]<=8'd241;
		data_a[18148]<=8'd248;
		data_a[18149]<=8'd249;
		data_a[18150]<=8'd255;
		data_a[18151]<=8'd99;
		data_a[18152]<=8'd84;
		data_a[18153]<=8'd85;
		data_a[18154]<=8'd88;
		data_a[18155]<=8'd83;
		data_a[18156]<=8'd74;
		data_a[18157]<=8'd69;
		data_a[18158]<=8'd53;
		data_a[18159]<=8'd83;
		data_a[18160]<=8'd73;
		data_a[18161]<=8'd77;
		data_a[18162]<=8'd78;
		data_a[18163]<=8'd79;
		data_a[18164]<=8'd68;
		data_a[18165]<=8'd76;
		data_a[18166]<=8'd73;
		data_a[18167]<=8'd75;
		data_a[18168]<=8'd63;
		data_a[18169]<=8'd65;
		data_a[18170]<=8'd61;
		data_a[18171]<=8'd161;
		data_a[18172]<=8'd164;
		data_a[18173]<=8'd169;
		data_a[18174]<=8'd174;
		data_a[18175]<=8'd175;
		data_a[18176]<=8'd171;
		data_a[18177]<=8'd180;
		data_a[18178]<=8'd185;
		data_a[18179]<=8'd192;
		data_a[18180]<=8'd159;
		data_a[18181]<=8'd90;
		data_a[18182]<=8'd99;
		data_a[18183]<=8'd103;
		data_a[18184]<=8'd104;
		data_a[18185]<=8'd109;
		data_a[18186]<=8'd103;
		data_a[18187]<=8'd111;
		data_a[18188]<=8'd118;
		data_a[18189]<=8'd115;
		data_a[18190]<=8'd114;
		data_a[18191]<=8'd113;
		data_a[18192]<=8'd104;
		data_a[18193]<=8'd100;
		data_a[18194]<=8'd101;
		data_a[18195]<=8'd97;
		data_a[18196]<=8'd100;
		data_a[18197]<=8'd104;
		data_a[18198]<=8'd101;
		data_a[18199]<=8'd94;
		data_a[18200]<=8'd94;
		data_a[18201]<=8'd100;
		data_a[18202]<=8'd102;
		data_a[18203]<=8'd95;
		data_a[18204]<=8'd100;
		data_a[18205]<=8'd94;
		data_a[18206]<=8'd99;
		data_a[18207]<=8'd107;
		data_a[18208]<=8'd108;
		data_a[18209]<=8'd103;
		data_a[18210]<=8'd125;
		data_a[18211]<=8'd223;
		data_a[18212]<=8'd231;
		data_a[18213]<=8'd232;
		data_a[18214]<=8'd232;
		data_a[18215]<=8'd234;
		data_a[18216]<=8'd236;
		data_a[18217]<=8'd235;
		data_a[18218]<=8'd234;
		data_a[18219]<=8'd234;
		data_a[18220]<=8'd235;
		data_a[18221]<=8'd237;
		data_a[18222]<=8'd235;
		data_a[18223]<=8'd235;
		data_a[18224]<=8'd234;
		data_a[18225]<=8'd234;
		data_a[18226]<=8'd237;
		data_a[18227]<=8'd242;
		data_a[18228]<=8'd244;
		data_a[18229]<=8'd242;
		data_a[18230]<=8'd240;
		data_a[18231]<=8'd245;
		data_a[18232]<=8'd243;
		data_a[18233]<=8'd243;
		data_a[18234]<=8'd241;
		data_a[18235]<=8'd246;
		data_a[18236]<=8'd244;
		data_a[18237]<=8'd241;
		data_a[18238]<=8'd243;
		data_a[18239]<=8'd175;
		data_a[18240]<=8'd60;
		data_a[18241]<=8'd65;
		data_a[18242]<=8'd66;
		data_a[18243]<=8'd58;
		data_a[18244]<=8'd68;
		data_a[18245]<=8'd82;
		data_a[18246]<=8'd84;
		data_a[18247]<=8'd89;
		data_a[18248]<=8'd111;
		data_a[18249]<=8'd107;
		data_a[18250]<=8'd112;
		data_a[18251]<=8'd117;
		data_a[18252]<=8'd114;
		data_a[18253]<=8'd118;
		data_a[18254]<=8'd112;
		data_a[18255]<=8'd113;
		data_a[18256]<=8'd111;
		data_a[18257]<=8'd108;
		data_a[18258]<=8'd110;
		data_a[18259]<=8'd94;
		data_a[18260]<=8'd91;
		data_a[18261]<=8'd92;
		data_a[18262]<=8'd89;
		data_a[18263]<=8'd90;
		data_a[18264]<=8'd82;
		data_a[18265]<=8'd83;
		data_a[18266]<=8'd79;
		data_a[18267]<=8'd76;
		data_a[18268]<=8'd63;
		data_a[18269]<=8'd61;
		data_a[18270]<=8'd50;
		data_a[18271]<=8'd54;
		data_a[18272]<=8'd59;
		data_a[18273]<=8'd57;
		data_a[18274]<=8'd50;
		data_a[18275]<=8'd47;
		data_a[18276]<=8'd49;
		data_a[18277]<=8'd50;
		data_a[18278]<=8'd72;
		data_a[18279]<=8'd78;
		data_a[18280]<=8'd109;
		data_a[18281]<=8'd149;
		data_a[18282]<=8'd147;
		data_a[18283]<=8'd145;
		data_a[18284]<=8'd66;
		data_a[18285]<=8'd68;
		data_a[18286]<=8'd77;
		data_a[18287]<=8'd95;
		data_a[18288]<=8'd113;
		data_a[18289]<=8'd121;
		data_a[18290]<=8'd131;
		data_a[18291]<=8'd247;
		data_a[18292]<=8'd244;
		data_a[18293]<=8'd243;
		data_a[18294]<=8'd249;
		data_a[18295]<=8'd241;
		data_a[18296]<=8'd241;
		data_a[18297]<=8'd246;
		data_a[18298]<=8'd245;
		data_a[18299]<=8'd244;
		data_a[18300]<=8'd255;
		data_a[18301]<=8'd58;
		data_a[18302]<=8'd58;
		data_a[18303]<=8'd71;
		data_a[18304]<=8'd78;
		data_a[18305]<=8'd78;
		data_a[18306]<=8'd70;
		data_a[18307]<=8'd72;
		data_a[18308]<=8'd52;
		data_a[18309]<=8'd74;
		data_a[18310]<=8'd73;
		data_a[18311]<=8'd74;
		data_a[18312]<=8'd75;
		data_a[18313]<=8'd76;
		data_a[18314]<=8'd76;
		data_a[18315]<=8'd78;
		data_a[18316]<=8'd74;
		data_a[18317]<=8'd68;
		data_a[18318]<=8'd68;
		data_a[18319]<=8'd59;
		data_a[18320]<=8'd71;
		data_a[18321]<=8'd161;
		data_a[18322]<=8'd163;
		data_a[18323]<=8'd168;
		data_a[18324]<=8'd167;
		data_a[18325]<=8'd173;
		data_a[18326]<=8'd178;
		data_a[18327]<=8'd188;
		data_a[18328]<=8'd187;
		data_a[18329]<=8'd187;
		data_a[18330]<=8'd181;
		data_a[18331]<=8'd75;
		data_a[18332]<=8'd92;
		data_a[18333]<=8'd99;
		data_a[18334]<=8'd101;
		data_a[18335]<=8'd103;
		data_a[18336]<=8'd101;
		data_a[18337]<=8'd108;
		data_a[18338]<=8'd116;
		data_a[18339]<=8'd115;
		data_a[18340]<=8'd117;
		data_a[18341]<=8'd109;
		data_a[18342]<=8'd108;
		data_a[18343]<=8'd96;
		data_a[18344]<=8'd91;
		data_a[18345]<=8'd86;
		data_a[18346]<=8'd88;
		data_a[18347]<=8'd91;
		data_a[18348]<=8'd87;
		data_a[18349]<=8'd87;
		data_a[18350]<=8'd95;
		data_a[18351]<=8'd107;
		data_a[18352]<=8'd101;
		data_a[18353]<=8'd95;
		data_a[18354]<=8'd104;
		data_a[18355]<=8'd90;
		data_a[18356]<=8'd96;
		data_a[18357]<=8'd102;
		data_a[18358]<=8'd102;
		data_a[18359]<=8'd120;
		data_a[18360]<=8'd163;
		data_a[18361]<=8'd241;
		data_a[18362]<=8'd229;
		data_a[18363]<=8'd235;
		data_a[18364]<=8'd233;
		data_a[18365]<=8'd234;
		data_a[18366]<=8'd235;
		data_a[18367]<=8'd235;
		data_a[18368]<=8'd235;
		data_a[18369]<=8'd235;
		data_a[18370]<=8'd236;
		data_a[18371]<=8'd237;
		data_a[18372]<=8'd235;
		data_a[18373]<=8'd236;
		data_a[18374]<=8'd235;
		data_a[18375]<=8'd234;
		data_a[18376]<=8'd237;
		data_a[18377]<=8'd242;
		data_a[18378]<=8'd243;
		data_a[18379]<=8'd241;
		data_a[18380]<=8'd241;
		data_a[18381]<=8'd242;
		data_a[18382]<=8'd241;
		data_a[18383]<=8'd245;
		data_a[18384]<=8'd242;
		data_a[18385]<=8'd242;
		data_a[18386]<=8'd240;
		data_a[18387]<=8'd241;
		data_a[18388]<=8'd249;
		data_a[18389]<=8'd207;
		data_a[18390]<=8'd91;
		data_a[18391]<=8'd70;
		data_a[18392]<=8'd62;
		data_a[18393]<=8'd69;
		data_a[18394]<=8'd61;
		data_a[18395]<=8'd71;
		data_a[18396]<=8'd75;
		data_a[18397]<=8'd81;
		data_a[18398]<=8'd102;
		data_a[18399]<=8'd103;
		data_a[18400]<=8'd100;
		data_a[18401]<=8'd112;
		data_a[18402]<=8'd102;
		data_a[18403]<=8'd112;
		data_a[18404]<=8'd111;
		data_a[18405]<=8'd105;
		data_a[18406]<=8'd107;
		data_a[18407]<=8'd103;
		data_a[18408]<=8'd104;
		data_a[18409]<=8'd88;
		data_a[18410]<=8'd91;
		data_a[18411]<=8'd90;
		data_a[18412]<=8'd79;
		data_a[18413]<=8'd75;
		data_a[18414]<=8'd75;
		data_a[18415]<=8'd79;
		data_a[18416]<=8'd65;
		data_a[18417]<=8'd69;
		data_a[18418]<=8'd58;
		data_a[18419]<=8'd55;
		data_a[18420]<=8'd53;
		data_a[18421]<=8'd50;
		data_a[18422]<=8'd60;
		data_a[18423]<=8'd54;
		data_a[18424]<=8'd42;
		data_a[18425]<=8'd48;
		data_a[18426]<=8'd52;
		data_a[18427]<=8'd54;
		data_a[18428]<=8'd73;
		data_a[18429]<=8'd101;
		data_a[18430]<=8'd117;
		data_a[18431]<=8'd150;
		data_a[18432]<=8'd145;
		data_a[18433]<=8'd140;
		data_a[18434]<=8'd83;
		data_a[18435]<=8'd62;
		data_a[18436]<=8'd80;
		data_a[18437]<=8'd87;
		data_a[18438]<=8'd98;
		data_a[18439]<=8'd114;
		data_a[18440]<=8'd136;
		data_a[18441]<=8'd244;
		data_a[18442]<=8'd240;
		data_a[18443]<=8'd241;
		data_a[18444]<=8'd240;
		data_a[18445]<=8'd241;
		data_a[18446]<=8'd250;
		data_a[18447]<=8'd242;
		data_a[18448]<=8'd142;
		data_a[18449]<=8'd124;
		data_a[18450]<=8'd254;
		data_a[18451]<=8'd74;
		data_a[18452]<=8'd70;
		data_a[18453]<=8'd72;
		data_a[18454]<=8'd75;
		data_a[18455]<=8'd59;
		data_a[18456]<=8'd57;
		data_a[18457]<=8'd60;
		data_a[18458]<=8'd59;
		data_a[18459]<=8'd57;
		data_a[18460]<=8'd82;
		data_a[18461]<=8'd76;
		data_a[18462]<=8'd76;
		data_a[18463]<=8'd73;
		data_a[18464]<=8'd74;
		data_a[18465]<=8'd67;
		data_a[18466]<=8'd72;
		data_a[18467]<=8'd67;
		data_a[18468]<=8'd56;
		data_a[18469]<=8'd62;
		data_a[18470]<=8'd68;
		data_a[18471]<=8'd156;
		data_a[18472]<=8'd172;
		data_a[18473]<=8'd163;
		data_a[18474]<=8'd176;
		data_a[18475]<=8'd172;
		data_a[18476]<=8'd177;
		data_a[18477]<=8'd180;
		data_a[18478]<=8'd182;
		data_a[18479]<=8'd189;
		data_a[18480]<=8'd189;
		data_a[18481]<=8'd82;
		data_a[18482]<=8'd84;
		data_a[18483]<=8'd93;
		data_a[18484]<=8'd96;
		data_a[18485]<=8'd98;
		data_a[18486]<=8'd98;
		data_a[18487]<=8'd104;
		data_a[18488]<=8'd114;
		data_a[18489]<=8'd117;
		data_a[18490]<=8'd113;
		data_a[18491]<=8'd106;
		data_a[18492]<=8'd104;
		data_a[18493]<=8'd97;
		data_a[18494]<=8'd93;
		data_a[18495]<=8'd85;
		data_a[18496]<=8'd78;
		data_a[18497]<=8'd74;
		data_a[18498]<=8'd83;
		data_a[18499]<=8'd84;
		data_a[18500]<=8'd92;
		data_a[18501]<=8'd98;
		data_a[18502]<=8'd90;
		data_a[18503]<=8'd91;
		data_a[18504]<=8'd100;
		data_a[18505]<=8'd91;
		data_a[18506]<=8'd99;
		data_a[18507]<=8'd107;
		data_a[18508]<=8'd111;
		data_a[18509]<=8'd118;
		data_a[18510]<=8'd201;
		data_a[18511]<=8'd224;
		data_a[18512]<=8'd237;
		data_a[18513]<=8'd232;
		data_a[18514]<=8'd234;
		data_a[18515]<=8'd234;
		data_a[18516]<=8'd235;
		data_a[18517]<=8'd235;
		data_a[18518]<=8'd235;
		data_a[18519]<=8'd235;
		data_a[18520]<=8'd236;
		data_a[18521]<=8'd236;
		data_a[18522]<=8'd235;
		data_a[18523]<=8'd236;
		data_a[18524]<=8'd235;
		data_a[18525]<=8'd234;
		data_a[18526]<=8'd237;
		data_a[18527]<=8'd242;
		data_a[18528]<=8'd244;
		data_a[18529]<=8'd241;
		data_a[18530]<=8'd243;
		data_a[18531]<=8'd242;
		data_a[18532]<=8'd242;
		data_a[18533]<=8'd247;
		data_a[18534]<=8'd243;
		data_a[18535]<=8'd240;
		data_a[18536]<=8'd237;
		data_a[18537]<=8'd241;
		data_a[18538]<=8'd244;
		data_a[18539]<=8'd210;
		data_a[18540]<=8'd136;
		data_a[18541]<=8'd65;
		data_a[18542]<=8'd61;
		data_a[18543]<=8'd60;
		data_a[18544]<=8'd67;
		data_a[18545]<=8'd70;
		data_a[18546]<=8'd70;
		data_a[18547]<=8'd81;
		data_a[18548]<=8'd88;
		data_a[18549]<=8'd98;
		data_a[18550]<=8'd99;
		data_a[18551]<=8'd105;
		data_a[18552]<=8'd105;
		data_a[18553]<=8'd106;
		data_a[18554]<=8'd100;
		data_a[18555]<=8'd97;
		data_a[18556]<=8'd85;
		data_a[18557]<=8'd89;
		data_a[18558]<=8'd92;
		data_a[18559]<=8'd78;
		data_a[18560]<=8'd73;
		data_a[18561]<=8'd86;
		data_a[18562]<=8'd72;
		data_a[18563]<=8'd72;
		data_a[18564]<=8'd70;
		data_a[18565]<=8'd64;
		data_a[18566]<=8'd63;
		data_a[18567]<=8'd62;
		data_a[18568]<=8'd47;
		data_a[18569]<=8'd54;
		data_a[18570]<=8'd46;
		data_a[18571]<=8'd47;
		data_a[18572]<=8'd56;
		data_a[18573]<=8'd55;
		data_a[18574]<=8'd46;
		data_a[18575]<=8'd52;
		data_a[18576]<=8'd52;
		data_a[18577]<=8'd56;
		data_a[18578]<=8'd78;
		data_a[18579]<=8'd103;
		data_a[18580]<=8'd135;
		data_a[18581]<=8'd141;
		data_a[18582]<=8'd144;
		data_a[18583]<=8'd142;
		data_a[18584]<=8'd92;
		data_a[18585]<=8'd60;
		data_a[18586]<=8'd73;
		data_a[18587]<=8'd84;
		data_a[18588]<=8'd94;
		data_a[18589]<=8'd115;
		data_a[18590]<=8'd127;
		data_a[18591]<=8'd245;
		data_a[18592]<=8'd249;
		data_a[18593]<=8'd238;
		data_a[18594]<=8'd245;
		data_a[18595]<=8'd248;
		data_a[18596]<=8'd164;
		data_a[18597]<=8'd133;
		data_a[18598]<=8'd142;
		data_a[18599]<=8'd146;
		data_a[18600]<=8'd255;
		data_a[18601]<=8'd51;
		data_a[18602]<=8'd65;
		data_a[18603]<=8'd62;
		data_a[18604]<=8'd63;
		data_a[18605]<=8'd71;
		data_a[18606]<=8'd70;
		data_a[18607]<=8'd69;
		data_a[18608]<=8'd64;
		data_a[18609]<=8'd65;
		data_a[18610]<=8'd75;
		data_a[18611]<=8'd75;
		data_a[18612]<=8'd76;
		data_a[18613]<=8'd79;
		data_a[18614]<=8'd71;
		data_a[18615]<=8'd79;
		data_a[18616]<=8'd71;
		data_a[18617]<=8'd65;
		data_a[18618]<=8'd55;
		data_a[18619]<=8'd61;
		data_a[18620]<=8'd52;
		data_a[18621]<=8'd161;
		data_a[18622]<=8'd165;
		data_a[18623]<=8'd175;
		data_a[18624]<=8'd172;
		data_a[18625]<=8'd173;
		data_a[18626]<=8'd178;
		data_a[18627]<=8'd183;
		data_a[18628]<=8'd189;
		data_a[18629]<=8'd193;
		data_a[18630]<=8'd189;
		data_a[18631]<=8'd110;
		data_a[18632]<=8'd80;
		data_a[18633]<=8'd88;
		data_a[18634]<=8'd93;
		data_a[18635]<=8'd97;
		data_a[18636]<=8'd99;
		data_a[18637]<=8'd103;
		data_a[18638]<=8'd114;
		data_a[18639]<=8'd118;
		data_a[18640]<=8'd122;
		data_a[18641]<=8'd117;
		data_a[18642]<=8'd99;
		data_a[18643]<=8'd93;
		data_a[18644]<=8'd90;
		data_a[18645]<=8'd89;
		data_a[18646]<=8'd87;
		data_a[18647]<=8'd89;
		data_a[18648]<=8'd86;
		data_a[18649]<=8'd89;
		data_a[18650]<=8'd97;
		data_a[18651]<=8'd96;
		data_a[18652]<=8'd94;
		data_a[18653]<=8'd98;
		data_a[18654]<=8'd95;
		data_a[18655]<=8'd96;
		data_a[18656]<=8'd95;
		data_a[18657]<=8'd105;
		data_a[18658]<=8'd102;
		data_a[18659]<=8'd87;
		data_a[18660]<=8'd236;
		data_a[18661]<=8'd231;
		data_a[18662]<=8'd233;
		data_a[18663]<=8'd233;
		data_a[18664]<=8'd234;
		data_a[18665]<=8'd234;
		data_a[18666]<=8'd234;
		data_a[18667]<=8'd235;
		data_a[18668]<=8'd235;
		data_a[18669]<=8'd236;
		data_a[18670]<=8'd236;
		data_a[18671]<=8'd236;
		data_a[18672]<=8'd235;
		data_a[18673]<=8'd236;
		data_a[18674]<=8'd234;
		data_a[18675]<=8'd233;
		data_a[18676]<=8'd237;
		data_a[18677]<=8'd242;
		data_a[18678]<=8'd244;
		data_a[18679]<=8'd242;
		data_a[18680]<=8'd241;
		data_a[18681]<=8'd246;
		data_a[18682]<=8'd245;
		data_a[18683]<=8'd244;
		data_a[18684]<=8'd240;
		data_a[18685]<=8'd244;
		data_a[18686]<=8'd241;
		data_a[18687]<=8'd239;
		data_a[18688]<=8'd248;
		data_a[18689]<=8'd241;
		data_a[18690]<=8'd131;
		data_a[18691]<=8'd70;
		data_a[18692]<=8'd63;
		data_a[18693]<=8'd60;
		data_a[18694]<=8'd70;
		data_a[18695]<=8'd62;
		data_a[18696]<=8'd67;
		data_a[18697]<=8'd74;
		data_a[18698]<=8'd82;
		data_a[18699]<=8'd83;
		data_a[18700]<=8'd96;
		data_a[18701]<=8'd85;
		data_a[18702]<=8'd100;
		data_a[18703]<=8'd91;
		data_a[18704]<=8'd96;
		data_a[18705]<=8'd84;
		data_a[18706]<=8'd80;
		data_a[18707]<=8'd91;
		data_a[18708]<=8'd73;
		data_a[18709]<=8'd68;
		data_a[18710]<=8'd72;
		data_a[18711]<=8'd74;
		data_a[18712]<=8'd69;
		data_a[18713]<=8'd61;
		data_a[18714]<=8'd66;
		data_a[18715]<=8'd65;
		data_a[18716]<=8'd56;
		data_a[18717]<=8'd62;
		data_a[18718]<=8'd54;
		data_a[18719]<=8'd52;
		data_a[18720]<=8'd52;
		data_a[18721]<=8'd54;
		data_a[18722]<=8'd46;
		data_a[18723]<=8'd44;
		data_a[18724]<=8'd42;
		data_a[18725]<=8'd48;
		data_a[18726]<=8'd53;
		data_a[18727]<=8'd67;
		data_a[18728]<=8'd97;
		data_a[18729]<=8'd104;
		data_a[18730]<=8'd132;
		data_a[18731]<=8'd141;
		data_a[18732]<=8'd144;
		data_a[18733]<=8'd134;
		data_a[18734]<=8'd108;
		data_a[18735]<=8'd56;
		data_a[18736]<=8'd73;
		data_a[18737]<=8'd81;
		data_a[18738]<=8'd95;
		data_a[18739]<=8'd96;
		data_a[18740]<=8'd121;
		data_a[18741]<=8'd228;
		data_a[18742]<=8'd244;
		data_a[18743]<=8'd228;
		data_a[18744]<=8'd152;
		data_a[18745]<=8'd130;
		data_a[18746]<=8'd127;
		data_a[18747]<=8'd130;
		data_a[18748]<=8'd125;
		data_a[18749]<=8'd122;
		data_a[18750]<=8'd255;
		data_a[18751]<=8'd66;
		data_a[18752]<=8'd59;
		data_a[18753]<=8'd55;
		data_a[18754]<=8'd54;
		data_a[18755]<=8'd44;
		data_a[18756]<=8'd48;
		data_a[18757]<=8'd53;
		data_a[18758]<=8'd61;
		data_a[18759]<=8'd67;
		data_a[18760]<=8'd63;
		data_a[18761]<=8'd67;
		data_a[18762]<=8'd67;
		data_a[18763]<=8'd68;
		data_a[18764]<=8'd64;
		data_a[18765]<=8'd73;
		data_a[18766]<=8'd73;
		data_a[18767]<=8'd67;
		data_a[18768]<=8'd43;
		data_a[18769]<=8'd52;
		data_a[18770]<=8'd66;
		data_a[18771]<=8'd167;
		data_a[18772]<=8'd170;
		data_a[18773]<=8'd166;
		data_a[18774]<=8'd170;
		data_a[18775]<=8'd179;
		data_a[18776]<=8'd176;
		data_a[18777]<=8'd183;
		data_a[18778]<=8'd187;
		data_a[18779]<=8'd186;
		data_a[18780]<=8'd191;
		data_a[18781]<=8'd147;
		data_a[18782]<=8'd77;
		data_a[18783]<=8'd79;
		data_a[18784]<=8'd86;
		data_a[18785]<=8'd93;
		data_a[18786]<=8'd98;
		data_a[18787]<=8'd100;
		data_a[18788]<=8'd114;
		data_a[18789]<=8'd118;
		data_a[18790]<=8'd111;
		data_a[18791]<=8'd115;
		data_a[18792]<=8'd101;
		data_a[18793]<=8'd97;
		data_a[18794]<=8'd90;
		data_a[18795]<=8'd84;
		data_a[18796]<=8'd79;
		data_a[18797]<=8'd81;
		data_a[18798]<=8'd78;
		data_a[18799]<=8'd82;
		data_a[18800]<=8'd92;
		data_a[18801]<=8'd93;
		data_a[18802]<=8'd96;
		data_a[18803]<=8'd99;
		data_a[18804]<=8'd86;
		data_a[18805]<=8'd91;
		data_a[18806]<=8'd105;
		data_a[18807]<=8'd104;
		data_a[18808]<=8'd108;
		data_a[18809]<=8'd168;
		data_a[18810]<=8'd238;
		data_a[18811]<=8'd237;
		data_a[18812]<=8'd231;
		data_a[18813]<=8'd237;
		data_a[18814]<=8'd234;
		data_a[18815]<=8'd234;
		data_a[18816]<=8'd235;
		data_a[18817]<=8'd235;
		data_a[18818]<=8'd235;
		data_a[18819]<=8'd236;
		data_a[18820]<=8'd236;
		data_a[18821]<=8'd236;
		data_a[18822]<=8'd236;
		data_a[18823]<=8'd236;
		data_a[18824]<=8'd234;
		data_a[18825]<=8'd233;
		data_a[18826]<=8'd236;
		data_a[18827]<=8'd242;
		data_a[18828]<=8'd245;
		data_a[18829]<=8'd243;
		data_a[18830]<=8'd242;
		data_a[18831]<=8'd244;
		data_a[18832]<=8'd243;
		data_a[18833]<=8'd245;
		data_a[18834]<=8'd242;
		data_a[18835]<=8'd244;
		data_a[18836]<=8'd242;
		data_a[18837]<=8'd243;
		data_a[18838]<=8'd248;
		data_a[18839]<=8'd247;
		data_a[18840]<=8'd185;
		data_a[18841]<=8'd67;
		data_a[18842]<=8'd61;
		data_a[18843]<=8'd59;
		data_a[18844]<=8'd62;
		data_a[18845]<=8'd64;
		data_a[18846]<=8'd63;
		data_a[18847]<=8'd68;
		data_a[18848]<=8'd76;
		data_a[18849]<=8'd75;
		data_a[18850]<=8'd82;
		data_a[18851]<=8'd77;
		data_a[18852]<=8'd85;
		data_a[18853]<=8'd82;
		data_a[18854]<=8'd79;
		data_a[18855]<=8'd76;
		data_a[18856]<=8'd70;
		data_a[18857]<=8'd70;
		data_a[18858]<=8'd68;
		data_a[18859]<=8'd62;
		data_a[18860]<=8'd60;
		data_a[18861]<=8'd59;
		data_a[18862]<=8'd57;
		data_a[18863]<=8'd61;
		data_a[18864]<=8'd56;
		data_a[18865]<=8'd61;
		data_a[18866]<=8'd60;
		data_a[18867]<=8'd65;
		data_a[18868]<=8'd48;
		data_a[18869]<=8'd52;
		data_a[18870]<=8'd46;
		data_a[18871]<=8'd53;
		data_a[18872]<=8'd42;
		data_a[18873]<=8'd45;
		data_a[18874]<=8'd48;
		data_a[18875]<=8'd47;
		data_a[18876]<=8'd49;
		data_a[18877]<=8'd72;
		data_a[18878]<=8'd104;
		data_a[18879]<=8'd110;
		data_a[18880]<=8'd142;
		data_a[18881]<=8'd139;
		data_a[18882]<=8'd139;
		data_a[18883]<=8'd138;
		data_a[18884]<=8'd99;
		data_a[18885]<=8'd59;
		data_a[18886]<=8'd67;
		data_a[18887]<=8'd83;
		data_a[18888]<=8'd84;
		data_a[18889]<=8'd110;
		data_a[18890]<=8'd127;
		data_a[18891]<=8'd167;
		data_a[18892]<=8'd155;
		data_a[18893]<=8'd116;
		data_a[18894]<=8'd121;
		data_a[18895]<=8'd105;
		data_a[18896]<=8'd114;
		data_a[18897]<=8'd120;
		data_a[18898]<=8'd115;
		data_a[18899]<=8'd124;
		data_a[18900]<=8'd255;
		data_a[18901]<=8'd65;
		data_a[18902]<=8'd69;
		data_a[18903]<=8'd62;
		data_a[18904]<=8'd58;
		data_a[18905]<=8'd62;
		data_a[18906]<=8'd52;
		data_a[18907]<=8'd33;
		data_a[18908]<=8'd33;
		data_a[18909]<=8'd40;
		data_a[18910]<=8'd56;
		data_a[18911]<=8'd61;
		data_a[18912]<=8'd63;
		data_a[18913]<=8'd61;
		data_a[18914]<=8'd63;
		data_a[18915]<=8'd61;
		data_a[18916]<=8'd60;
		data_a[18917]<=8'd59;
		data_a[18918]<=8'd65;
		data_a[18919]<=8'd58;
		data_a[18920]<=8'd64;
		data_a[18921]<=8'd161;
		data_a[18922]<=8'd165;
		data_a[18923]<=8'd172;
		data_a[18924]<=8'd170;
		data_a[18925]<=8'd175;
		data_a[18926]<=8'd175;
		data_a[18927]<=8'd187;
		data_a[18928]<=8'd193;
		data_a[18929]<=8'd191;
		data_a[18930]<=8'd191;
		data_a[18931]<=8'd157;
		data_a[18932]<=8'd80;
		data_a[18933]<=8'd72;
		data_a[18934]<=8'd76;
		data_a[18935]<=8'd84;
		data_a[18936]<=8'd90;
		data_a[18937]<=8'd93;
		data_a[18938]<=8'd110;
		data_a[18939]<=8'd114;
		data_a[18940]<=8'd119;
		data_a[18941]<=8'd117;
		data_a[18942]<=8'd114;
		data_a[18943]<=8'd104;
		data_a[18944]<=8'd93;
		data_a[18945]<=8'd88;
		data_a[18946]<=8'd85;
		data_a[18947]<=8'd87;
		data_a[18948]<=8'd86;
		data_a[18949]<=8'd86;
		data_a[18950]<=8'd88;
		data_a[18951]<=8'd92;
		data_a[18952]<=8'd95;
		data_a[18953]<=8'd98;
		data_a[18954]<=8'd89;
		data_a[18955]<=8'd95;
		data_a[18956]<=8'd92;
		data_a[18957]<=8'd104;
		data_a[18958]<=8'd115;
		data_a[18959]<=8'd230;
		data_a[18960]<=8'd235;
		data_a[18961]<=8'd232;
		data_a[18962]<=8'd235;
		data_a[18963]<=8'd235;
		data_a[18964]<=8'd234;
		data_a[18965]<=8'd235;
		data_a[18966]<=8'd235;
		data_a[18967]<=8'd235;
		data_a[18968]<=8'd235;
		data_a[18969]<=8'd236;
		data_a[18970]<=8'd236;
		data_a[18971]<=8'd236;
		data_a[18972]<=8'd236;
		data_a[18973]<=8'd236;
		data_a[18974]<=8'd235;
		data_a[18975]<=8'd234;
		data_a[18976]<=8'd237;
		data_a[18977]<=8'd242;
		data_a[18978]<=8'd244;
		data_a[18979]<=8'd242;
		data_a[18980]<=8'd245;
		data_a[18981]<=8'd242;
		data_a[18982]<=8'd240;
		data_a[18983]<=8'd246;
		data_a[18984]<=8'd244;
		data_a[18985]<=8'd243;
		data_a[18986]<=8'd242;
		data_a[18987]<=8'd246;
		data_a[18988]<=8'd242;
		data_a[18989]<=8'd252;
		data_a[18990]<=8'd209;
		data_a[18991]<=8'd81;
		data_a[18992]<=8'd66;
		data_a[18993]<=8'd59;
		data_a[18994]<=8'd70;
		data_a[18995]<=8'd58;
		data_a[18996]<=8'd63;
		data_a[18997]<=8'd69;
		data_a[18998]<=8'd70;
		data_a[18999]<=8'd78;
		data_a[19000]<=8'd75;
		data_a[19001]<=8'd82;
		data_a[19002]<=8'd77;
		data_a[19003]<=8'd79;
		data_a[19004]<=8'd72;
		data_a[19005]<=8'd65;
		data_a[19006]<=8'd63;
		data_a[19007]<=8'd62;
		data_a[19008]<=8'd62;
		data_a[19009]<=8'd58;
		data_a[19010]<=8'd59;
		data_a[19011]<=8'd48;
		data_a[19012]<=8'd52;
		data_a[19013]<=8'd51;
		data_a[19014]<=8'd52;
		data_a[19015]<=8'd60;
		data_a[19016]<=8'd56;
		data_a[19017]<=8'd59;
		data_a[19018]<=8'd51;
		data_a[19019]<=8'd45;
		data_a[19020]<=8'd47;
		data_a[19021]<=8'd49;
		data_a[19022]<=8'd41;
		data_a[19023]<=8'd43;
		data_a[19024]<=8'd43;
		data_a[19025]<=8'd45;
		data_a[19026]<=8'd48;
		data_a[19027]<=8'd85;
		data_a[19028]<=8'd102;
		data_a[19029]<=8'd127;
		data_a[19030]<=8'd141;
		data_a[19031]<=8'd140;
		data_a[19032]<=8'd139;
		data_a[19033]<=8'd130;
		data_a[19034]<=8'd99;
		data_a[19035]<=8'd63;
		data_a[19036]<=8'd74;
		data_a[19037]<=8'd78;
		data_a[19038]<=8'd83;
		data_a[19039]<=8'd96;
		data_a[19040]<=8'd113;
		data_a[19041]<=8'd136;
		data_a[19042]<=8'd149;
		data_a[19043]<=8'd122;
		data_a[19044]<=8'd108;
		data_a[19045]<=8'd90;
		data_a[19046]<=8'd115;
		data_a[19047]<=8'd107;
		data_a[19048]<=8'd112;
		data_a[19049]<=8'd113;
		data_a[19050]<=8'd255;
		data_a[19051]<=8'd72;
		data_a[19052]<=8'd68;
		data_a[19053]<=8'd69;
		data_a[19054]<=8'd67;
		data_a[19055]<=8'd62;
		data_a[19056]<=8'd57;
		data_a[19057]<=8'd48;
		data_a[19058]<=8'd50;
		data_a[19059]<=8'd53;
		data_a[19060]<=8'd72;
		data_a[19061]<=8'd63;
		data_a[19062]<=8'd55;
		data_a[19063]<=8'd60;
		data_a[19064]<=8'd51;
		data_a[19065]<=8'd54;
		data_a[19066]<=8'd59;
		data_a[19067]<=8'd58;
		data_a[19068]<=8'd60;
		data_a[19069]<=8'd70;
		data_a[19070]<=8'd53;
		data_a[19071]<=8'd164;
		data_a[19072]<=8'd168;
		data_a[19073]<=8'd169;
		data_a[19074]<=8'd177;
		data_a[19075]<=8'd174;
		data_a[19076]<=8'd183;
		data_a[19077]<=8'd185;
		data_a[19078]<=8'd185;
		data_a[19079]<=8'd192;
		data_a[19080]<=8'd194;
		data_a[19081]<=8'd175;
		data_a[19082]<=8'd89;
		data_a[19083]<=8'd72;
		data_a[19084]<=8'd71;
		data_a[19085]<=8'd77;
		data_a[19086]<=8'd82;
		data_a[19087]<=8'd86;
		data_a[19088]<=8'd104;
		data_a[19089]<=8'd108;
		data_a[19090]<=8'd119;
		data_a[19091]<=8'd109;
		data_a[19092]<=8'd119;
		data_a[19093]<=8'd106;
		data_a[19094]<=8'd96;
		data_a[19095]<=8'd95;
		data_a[19096]<=8'd92;
		data_a[19097]<=8'd92;
		data_a[19098]<=8'd90;
		data_a[19099]<=8'd90;
		data_a[19100]<=8'd88;
		data_a[19101]<=8'd98;
		data_a[19102]<=8'd97;
		data_a[19103]<=8'd94;
		data_a[19104]<=8'd87;
		data_a[19105]<=8'd87;
		data_a[19106]<=8'd88;
		data_a[19107]<=8'd105;
		data_a[19108]<=8'd198;
		data_a[19109]<=8'd238;
		data_a[19110]<=8'd237;
		data_a[19111]<=8'd235;
		data_a[19112]<=8'd237;
		data_a[19113]<=8'd235;
		data_a[19114]<=8'd234;
		data_a[19115]<=8'd235;
		data_a[19116]<=8'd235;
		data_a[19117]<=8'd235;
		data_a[19118]<=8'd235;
		data_a[19119]<=8'd235;
		data_a[19120]<=8'd236;
		data_a[19121]<=8'd236;
		data_a[19122]<=8'd235;
		data_a[19123]<=8'd236;
		data_a[19124]<=8'd235;
		data_a[19125]<=8'd234;
		data_a[19126]<=8'd238;
		data_a[19127]<=8'd242;
		data_a[19128]<=8'd243;
		data_a[19129]<=8'd241;
		data_a[19130]<=8'd243;
		data_a[19131]<=8'd245;
		data_a[19132]<=8'd242;
		data_a[19133]<=8'd242;
		data_a[19134]<=8'd240;
		data_a[19135]<=8'd245;
		data_a[19136]<=8'd244;
		data_a[19137]<=8'd243;
		data_a[19138]<=8'd244;
		data_a[19139]<=8'd240;
		data_a[19140]<=8'd223;
		data_a[19141]<=8'd86;
		data_a[19142]<=8'd72;
		data_a[19143]<=8'd61;
		data_a[19144]<=8'd58;
		data_a[19145]<=8'd69;
		data_a[19146]<=8'd62;
		data_a[19147]<=8'd65;
		data_a[19148]<=8'd62;
		data_a[19149]<=8'd72;
		data_a[19150]<=8'd74;
		data_a[19151]<=8'd77;
		data_a[19152]<=8'd74;
		data_a[19153]<=8'd68;
		data_a[19154]<=8'd66;
		data_a[19155]<=8'd67;
		data_a[19156]<=8'd60;
		data_a[19157]<=8'd59;
		data_a[19158]<=8'd60;
		data_a[19159]<=8'd50;
		data_a[19160]<=8'd47;
		data_a[19161]<=8'd51;
		data_a[19162]<=8'd48;
		data_a[19163]<=8'd48;
		data_a[19164]<=8'd51;
		data_a[19165]<=8'd53;
		data_a[19166]<=8'd61;
		data_a[19167]<=8'd54;
		data_a[19168]<=8'd52;
		data_a[19169]<=8'd44;
		data_a[19170]<=8'd45;
		data_a[19171]<=8'd43;
		data_a[19172]<=8'd45;
		data_a[19173]<=8'd47;
		data_a[19174]<=8'd43;
		data_a[19175]<=8'd45;
		data_a[19176]<=8'd43;
		data_a[19177]<=8'd87;
		data_a[19178]<=8'd115;
		data_a[19179]<=8'd121;
		data_a[19180]<=8'd134;
		data_a[19181]<=8'd139;
		data_a[19182]<=8'd137;
		data_a[19183]<=8'd124;
		data_a[19184]<=8'd102;
		data_a[19185]<=8'd69;
		data_a[19186]<=8'd65;
		data_a[19187]<=8'd79;
		data_a[19188]<=8'd89;
		data_a[19189]<=8'd98;
		data_a[19190]<=8'd107;
		data_a[19191]<=8'd139;
		data_a[19192]<=8'd90;
		data_a[19193]<=8'd114;
		data_a[19194]<=8'd106;
		data_a[19195]<=8'd111;
		data_a[19196]<=8'd106;
		data_a[19197]<=8'd111;
		data_a[19198]<=8'd109;
		data_a[19199]<=8'd111;
		data_a[19200]<=8'd254;
		data_a[19201]<=8'd56;
		data_a[19202]<=8'd59;
		data_a[19203]<=8'd70;
		data_a[19204]<=8'd73;
		data_a[19205]<=8'd68;
		data_a[19206]<=8'd63;
		data_a[19207]<=8'd54;
		data_a[19208]<=8'd46;
		data_a[19209]<=8'd58;
		data_a[19210]<=8'd81;
		data_a[19211]<=8'd75;
		data_a[19212]<=8'd69;
		data_a[19213]<=8'd74;
		data_a[19214]<=8'd70;
		data_a[19215]<=8'd66;
		data_a[19216]<=8'd67;
		data_a[19217]<=8'd53;
		data_a[19218]<=8'd44;
		data_a[19219]<=8'd43;
		data_a[19220]<=8'd55;
		data_a[19221]<=8'd161;
		data_a[19222]<=8'd164;
		data_a[19223]<=8'd175;
		data_a[19224]<=8'd174;
		data_a[19225]<=8'd176;
		data_a[19226]<=8'd177;
		data_a[19227]<=8'd188;
		data_a[19228]<=8'd189;
		data_a[19229]<=8'd194;
		data_a[19230]<=8'd197;
		data_a[19231]<=8'd182;
		data_a[19232]<=8'd122;
		data_a[19233]<=8'd73;
		data_a[19234]<=8'd64;
		data_a[19235]<=8'd68;
		data_a[19236]<=8'd73;
		data_a[19237]<=8'd77;
		data_a[19238]<=8'd96;
		data_a[19239]<=8'd108;
		data_a[19240]<=8'd114;
		data_a[19241]<=8'd117;
		data_a[19242]<=8'd114;
		data_a[19243]<=8'd112;
		data_a[19244]<=8'd103;
		data_a[19245]<=8'd101;
		data_a[19246]<=8'd97;
		data_a[19247]<=8'd96;
		data_a[19248]<=8'd88;
		data_a[19249]<=8'd92;
		data_a[19250]<=8'd79;
		data_a[19251]<=8'd100;
		data_a[19252]<=8'd87;
		data_a[19253]<=8'd82;
		data_a[19254]<=8'd86;
		data_a[19255]<=8'd81;
		data_a[19256]<=8'd86;
		data_a[19257]<=8'd81;
		data_a[19258]<=8'd241;
		data_a[19259]<=8'd239;
		data_a[19260]<=8'd231;
		data_a[19261]<=8'd240;
		data_a[19262]<=8'd234;
		data_a[19263]<=8'd235;
		data_a[19264]<=8'd235;
		data_a[19265]<=8'd235;
		data_a[19266]<=8'd236;
		data_a[19267]<=8'd237;
		data_a[19268]<=8'd236;
		data_a[19269]<=8'd235;
		data_a[19270]<=8'd235;
		data_a[19271]<=8'd236;
		data_a[19272]<=8'd236;
		data_a[19273]<=8'd234;
		data_a[19274]<=8'd237;
		data_a[19275]<=8'd234;
		data_a[19276]<=8'd238;
		data_a[19277]<=8'd238;
		data_a[19278]<=8'd244;
		data_a[19279]<=8'd242;
		data_a[19280]<=8'd240;
		data_a[19281]<=8'd242;
		data_a[19282]<=8'd243;
		data_a[19283]<=8'd243;
		data_a[19284]<=8'd243;
		data_a[19285]<=8'd244;
		data_a[19286]<=8'd244;
		data_a[19287]<=8'd243;
		data_a[19288]<=8'd244;
		data_a[19289]<=8'd239;
		data_a[19290]<=8'd250;
		data_a[19291]<=8'd139;
		data_a[19292]<=8'd55;
		data_a[19293]<=8'd58;
		data_a[19294]<=8'd64;
		data_a[19295]<=8'd65;
		data_a[19296]<=8'd62;
		data_a[19297]<=8'd59;
		data_a[19298]<=8'd54;
		data_a[19299]<=8'd70;
		data_a[19300]<=8'd63;
		data_a[19301]<=8'd58;
		data_a[19302]<=8'd65;
		data_a[19303]<=8'd67;
		data_a[19304]<=8'd58;
		data_a[19305]<=8'd60;
		data_a[19306]<=8'd56;
		data_a[19307]<=8'd49;
		data_a[19308]<=8'd48;
		data_a[19309]<=8'd46;
		data_a[19310]<=8'd42;
		data_a[19311]<=8'd43;
		data_a[19312]<=8'd45;
		data_a[19313]<=8'd50;
		data_a[19314]<=8'd48;
		data_a[19315]<=8'd50;
		data_a[19316]<=8'd48;
		data_a[19317]<=8'd50;
		data_a[19318]<=8'd43;
		data_a[19319]<=8'd40;
		data_a[19320]<=8'd44;
		data_a[19321]<=8'd39;
		data_a[19322]<=8'd41;
		data_a[19323]<=8'd44;
		data_a[19324]<=8'd42;
		data_a[19325]<=8'd50;
		data_a[19326]<=8'd58;
		data_a[19327]<=8'd91;
		data_a[19328]<=8'd119;
		data_a[19329]<=8'd130;
		data_a[19330]<=8'd135;
		data_a[19331]<=8'd136;
		data_a[19332]<=8'd138;
		data_a[19333]<=8'd124;
		data_a[19334]<=8'd105;
		data_a[19335]<=8'd68;
		data_a[19336]<=8'd67;
		data_a[19337]<=8'd86;
		data_a[19338]<=8'd84;
		data_a[19339]<=8'd92;
		data_a[19340]<=8'd107;
		data_a[19341]<=8'd120;
		data_a[19342]<=8'd121;
		data_a[19343]<=8'd120;
		data_a[19344]<=8'd117;
		data_a[19345]<=8'd118;
		data_a[19346]<=8'd102;
		data_a[19347]<=8'd104;
		data_a[19348]<=8'd102;
		data_a[19349]<=8'd98;
		data_a[19350]<=8'd254;
		data_a[19351]<=8'd96;
		data_a[19352]<=8'd102;
		data_a[19353]<=8'd79;
		data_a[19354]<=8'd64;
		data_a[19355]<=8'd60;
		data_a[19356]<=8'd60;
		data_a[19357]<=8'd53;
		data_a[19358]<=8'd54;
		data_a[19359]<=8'd55;
		data_a[19360]<=8'd68;
		data_a[19361]<=8'd78;
		data_a[19362]<=8'd74;
		data_a[19363]<=8'd77;
		data_a[19364]<=8'd75;
		data_a[19365]<=8'd73;
		data_a[19366]<=8'd71;
		data_a[19367]<=8'd63;
		data_a[19368]<=8'd83;
		data_a[19369]<=8'd64;
		data_a[19370]<=8'd57;
		data_a[19371]<=8'd164;
		data_a[19372]<=8'd176;
		data_a[19373]<=8'd164;
		data_a[19374]<=8'd173;
		data_a[19375]<=8'd170;
		data_a[19376]<=8'd188;
		data_a[19377]<=8'd188;
		data_a[19378]<=8'd189;
		data_a[19379]<=8'd193;
		data_a[19380]<=8'd197;
		data_a[19381]<=8'd191;
		data_a[19382]<=8'd132;
		data_a[19383]<=8'd96;
		data_a[19384]<=8'd67;
		data_a[19385]<=8'd69;
		data_a[19386]<=8'd64;
		data_a[19387]<=8'd73;
		data_a[19388]<=8'd86;
		data_a[19389]<=8'd101;
		data_a[19390]<=8'd113;
		data_a[19391]<=8'd107;
		data_a[19392]<=8'd110;
		data_a[19393]<=8'd105;
		data_a[19394]<=8'd102;
		data_a[19395]<=8'd103;
		data_a[19396]<=8'd97;
		data_a[19397]<=8'd94;
		data_a[19398]<=8'd87;
		data_a[19399]<=8'd91;
		data_a[19400]<=8'd94;
		data_a[19401]<=8'd94;
		data_a[19402]<=8'd89;
		data_a[19403]<=8'd85;
		data_a[19404]<=8'd75;
		data_a[19405]<=8'd79;
		data_a[19406]<=8'd87;
		data_a[19407]<=8'd123;
		data_a[19408]<=8'd240;
		data_a[19409]<=8'd233;
		data_a[19410]<=8'd233;
		data_a[19411]<=8'd232;
		data_a[19412]<=8'd236;
		data_a[19413]<=8'd238;
		data_a[19414]<=8'd235;
		data_a[19415]<=8'd235;
		data_a[19416]<=8'd236;
		data_a[19417]<=8'd236;
		data_a[19418]<=8'd236;
		data_a[19419]<=8'd235;
		data_a[19420]<=8'd235;
		data_a[19421]<=8'd236;
		data_a[19422]<=8'd235;
		data_a[19423]<=8'd234;
		data_a[19424]<=8'd237;
		data_a[19425]<=8'd235;
		data_a[19426]<=8'd238;
		data_a[19427]<=8'd239;
		data_a[19428]<=8'd243;
		data_a[19429]<=8'd240;
		data_a[19430]<=8'd242;
		data_a[19431]<=8'd243;
		data_a[19432]<=8'd243;
		data_a[19433]<=8'd242;
		data_a[19434]<=8'd242;
		data_a[19435]<=8'd242;
		data_a[19436]<=8'd243;
		data_a[19437]<=8'd242;
		data_a[19438]<=8'd241;
		data_a[19439]<=8'd247;
		data_a[19440]<=8'd237;
		data_a[19441]<=8'd150;
		data_a[19442]<=8'd133;
		data_a[19443]<=8'd90;
		data_a[19444]<=8'd68;
		data_a[19445]<=8'd60;
		data_a[19446]<=8'd57;
		data_a[19447]<=8'd62;
		data_a[19448]<=8'd53;
		data_a[19449]<=8'd64;
		data_a[19450]<=8'd61;
		data_a[19451]<=8'd58;
		data_a[19452]<=8'd57;
		data_a[19453]<=8'd55;
		data_a[19454]<=8'd56;
		data_a[19455]<=8'd54;
		data_a[19456]<=8'd45;
		data_a[19457]<=8'd45;
		data_a[19458]<=8'd45;
		data_a[19459]<=8'd40;
		data_a[19460]<=8'd40;
		data_a[19461]<=8'd37;
		data_a[19462]<=8'd49;
		data_a[19463]<=8'd38;
		data_a[19464]<=8'd36;
		data_a[19465]<=8'd49;
		data_a[19466]<=8'd50;
		data_a[19467]<=8'd39;
		data_a[19468]<=8'd37;
		data_a[19469]<=8'd51;
		data_a[19470]<=8'd37;
		data_a[19471]<=8'd43;
		data_a[19472]<=8'd45;
		data_a[19473]<=8'd42;
		data_a[19474]<=8'd49;
		data_a[19475]<=8'd41;
		data_a[19476]<=8'd63;
		data_a[19477]<=8'd103;
		data_a[19478]<=8'd122;
		data_a[19479]<=8'd128;
		data_a[19480]<=8'd133;
		data_a[19481]<=8'd135;
		data_a[19482]<=8'd134;
		data_a[19483]<=8'd120;
		data_a[19484]<=8'd103;
		data_a[19485]<=8'd69;
		data_a[19486]<=8'd66;
		data_a[19487]<=8'd76;
		data_a[19488]<=8'd85;
		data_a[19489]<=8'd89;
		data_a[19490]<=8'd110;
		data_a[19491]<=8'd121;
		data_a[19492]<=8'd133;
		data_a[19493]<=8'd124;
		data_a[19494]<=8'd111;
		data_a[19495]<=8'd111;
		data_a[19496]<=8'd99;
		data_a[19497]<=8'd104;
		data_a[19498]<=8'd100;
		data_a[19499]<=8'd95;
		data_a[19500]<=8'd254;
		data_a[19501]<=8'd94;
		data_a[19502]<=8'd99;
		data_a[19503]<=8'd90;
		data_a[19504]<=8'd84;
		data_a[19505]<=8'd65;
		data_a[19506]<=8'd55;
		data_a[19507]<=8'd57;
		data_a[19508]<=8'd50;
		data_a[19509]<=8'd65;
		data_a[19510]<=8'd81;
		data_a[19511]<=8'd77;
		data_a[19512]<=8'd75;
		data_a[19513]<=8'd77;
		data_a[19514]<=8'd70;
		data_a[19515]<=8'd72;
		data_a[19516]<=8'd87;
		data_a[19517]<=8'd121;
		data_a[19518]<=8'd109;
		data_a[19519]<=8'd129;
		data_a[19520]<=8'd101;
		data_a[19521]<=8'd159;
		data_a[19522]<=8'd173;
		data_a[19523]<=8'd174;
		data_a[19524]<=8'd174;
		data_a[19525]<=8'd180;
		data_a[19526]<=8'd175;
		data_a[19527]<=8'd188;
		data_a[19528]<=8'd196;
		data_a[19529]<=8'd195;
		data_a[19530]<=8'd192;
		data_a[19531]<=8'd197;
		data_a[19532]<=8'd139;
		data_a[19533]<=8'd113;
		data_a[19534]<=8'd67;
		data_a[19535]<=8'd62;
		data_a[19536]<=8'd63;
		data_a[19537]<=8'd73;
		data_a[19538]<=8'd81;
		data_a[19539]<=8'd92;
		data_a[19540]<=8'd106;
		data_a[19541]<=8'd95;
		data_a[19542]<=8'd105;
		data_a[19543]<=8'd99;
		data_a[19544]<=8'd100;
		data_a[19545]<=8'd103;
		data_a[19546]<=8'd100;
		data_a[19547]<=8'd96;
		data_a[19548]<=8'd93;
		data_a[19549]<=8'd94;
		data_a[19550]<=8'd93;
		data_a[19551]<=8'd90;
		data_a[19552]<=8'd78;
		data_a[19553]<=8'd75;
		data_a[19554]<=8'd79;
		data_a[19555]<=8'd74;
		data_a[19556]<=8'd80;
		data_a[19557]<=8'd141;
		data_a[19558]<=8'd235;
		data_a[19559]<=8'd234;
		data_a[19560]<=8'd240;
		data_a[19561]<=8'd232;
		data_a[19562]<=8'd234;
		data_a[19563]<=8'd233;
		data_a[19564]<=8'd235;
		data_a[19565]<=8'd235;
		data_a[19566]<=8'd235;
		data_a[19567]<=8'd236;
		data_a[19568]<=8'd236;
		data_a[19569]<=8'd235;
		data_a[19570]<=8'd235;
		data_a[19571]<=8'd236;
		data_a[19572]<=8'd235;
		data_a[19573]<=8'd234;
		data_a[19574]<=8'd237;
		data_a[19575]<=8'd236;
		data_a[19576]<=8'd238;
		data_a[19577]<=8'd239;
		data_a[19578]<=8'd242;
		data_a[19579]<=8'd239;
		data_a[19580]<=8'd243;
		data_a[19581]<=8'd243;
		data_a[19582]<=8'd243;
		data_a[19583]<=8'd241;
		data_a[19584]<=8'd241;
		data_a[19585]<=8'd241;
		data_a[19586]<=8'd242;
		data_a[19587]<=8'd242;
		data_a[19588]<=8'd241;
		data_a[19589]<=8'd247;
		data_a[19590]<=8'd235;
		data_a[19591]<=8'd250;
		data_a[19592]<=8'd225;
		data_a[19593]<=8'd164;
		data_a[19594]<=8'd59;
		data_a[19595]<=8'd69;
		data_a[19596]<=8'd62;
		data_a[19597]<=8'd59;
		data_a[19598]<=8'd54;
		data_a[19599]<=8'd49;
		data_a[19600]<=8'd50;
		data_a[19601]<=8'd54;
		data_a[19602]<=8'd41;
		data_a[19603]<=8'd56;
		data_a[19604]<=8'd52;
		data_a[19605]<=8'd48;
		data_a[19606]<=8'd51;
		data_a[19607]<=8'd43;
		data_a[19608]<=8'd37;
		data_a[19609]<=8'd39;
		data_a[19610]<=8'd36;
		data_a[19611]<=8'd39;
		data_a[19612]<=8'd38;
		data_a[19613]<=8'd45;
		data_a[19614]<=8'd44;
		data_a[19615]<=8'd35;
		data_a[19616]<=8'd38;
		data_a[19617]<=8'd43;
		data_a[19618]<=8'd45;
		data_a[19619]<=8'd41;
		data_a[19620]<=8'd45;
		data_a[19621]<=8'd47;
		data_a[19622]<=8'd33;
		data_a[19623]<=8'd38;
		data_a[19624]<=8'd43;
		data_a[19625]<=8'd46;
		data_a[19626]<=8'd77;
		data_a[19627]<=8'd112;
		data_a[19628]<=8'd126;
		data_a[19629]<=8'd127;
		data_a[19630]<=8'd131;
		data_a[19631]<=8'd134;
		data_a[19632]<=8'd129;
		data_a[19633]<=8'd116;
		data_a[19634]<=8'd101;
		data_a[19635]<=8'd70;
		data_a[19636]<=8'd74;
		data_a[19637]<=8'd78;
		data_a[19638]<=8'd84;
		data_a[19639]<=8'd92;
		data_a[19640]<=8'd99;
		data_a[19641]<=8'd118;
		data_a[19642]<=8'd126;
		data_a[19643]<=8'd114;
		data_a[19644]<=8'd104;
		data_a[19645]<=8'd102;
		data_a[19646]<=8'd96;
		data_a[19647]<=8'd103;
		data_a[19648]<=8'd98;
		data_a[19649]<=8'd91;
		data_a[19650]<=8'd253;
		data_a[19651]<=8'd89;
		data_a[19652]<=8'd91;
		data_a[19653]<=8'd85;
		data_a[19654]<=8'd84;
		data_a[19655]<=8'd66;
		data_a[19656]<=8'd56;
		data_a[19657]<=8'd57;
		data_a[19658]<=8'd51;
		data_a[19659]<=8'd62;
		data_a[19660]<=8'd74;
		data_a[19661]<=8'd72;
		data_a[19662]<=8'd77;
		data_a[19663]<=8'd67;
		data_a[19664]<=8'd83;
		data_a[19665]<=8'd109;
		data_a[19666]<=8'd92;
		data_a[19667]<=8'd93;
		data_a[19668]<=8'd84;
		data_a[19669]<=8'd144;
		data_a[19670]<=8'd73;
		data_a[19671]<=8'd160;
		data_a[19672]<=8'd165;
		data_a[19673]<=8'd172;
		data_a[19674]<=8'd178;
		data_a[19675]<=8'd177;
		data_a[19676]<=8'd186;
		data_a[19677]<=8'd187;
		data_a[19678]<=8'd192;
		data_a[19679]<=8'd197;
		data_a[19680]<=8'd199;
		data_a[19681]<=8'd185;
		data_a[19682]<=8'd136;
		data_a[19683]<=8'd127;
		data_a[19684]<=8'd91;
		data_a[19685]<=8'd61;
		data_a[19686]<=8'd62;
		data_a[19687]<=8'd59;
		data_a[19688]<=8'd70;
		data_a[19689]<=8'd86;
		data_a[19690]<=8'd95;
		data_a[19691]<=8'd88;
		data_a[19692]<=8'd98;
		data_a[19693]<=8'd98;
		data_a[19694]<=8'd96;
		data_a[19695]<=8'd102;
		data_a[19696]<=8'd105;
		data_a[19697]<=8'd100;
		data_a[19698]<=8'd93;
		data_a[19699]<=8'd94;
		data_a[19700]<=8'd87;
		data_a[19701]<=8'd91;
		data_a[19702]<=8'd74;
		data_a[19703]<=8'd73;
		data_a[19704]<=8'd73;
		data_a[19705]<=8'd73;
		data_a[19706]<=8'd105;
		data_a[19707]<=8'd142;
		data_a[19708]<=8'd236;
		data_a[19709]<=8'd235;
		data_a[19710]<=8'd236;
		data_a[19711]<=8'd235;
		data_a[19712]<=8'd234;
		data_a[19713]<=8'd235;
		data_a[19714]<=8'd235;
		data_a[19715]<=8'd235;
		data_a[19716]<=8'd235;
		data_a[19717]<=8'd236;
		data_a[19718]<=8'd236;
		data_a[19719]<=8'd235;
		data_a[19720]<=8'd235;
		data_a[19721]<=8'd236;
		data_a[19722]<=8'd236;
		data_a[19723]<=8'd234;
		data_a[19724]<=8'd235;
		data_a[19725]<=8'd235;
		data_a[19726]<=8'd236;
		data_a[19727]<=8'd239;
		data_a[19728]<=8'd242;
		data_a[19729]<=8'd240;
		data_a[19730]<=8'd242;
		data_a[19731]<=8'd242;
		data_a[19732]<=8'd242;
		data_a[19733]<=8'd241;
		data_a[19734]<=8'd241;
		data_a[19735]<=8'd241;
		data_a[19736]<=8'd241;
		data_a[19737]<=8'd242;
		data_a[19738]<=8'd245;
		data_a[19739]<=8'd233;
		data_a[19740]<=8'd239;
		data_a[19741]<=8'd227;
		data_a[19742]<=8'd246;
		data_a[19743]<=8'd242;
		data_a[19744]<=8'd109;
		data_a[19745]<=8'd67;
		data_a[19746]<=8'd61;
		data_a[19747]<=8'd55;
		data_a[19748]<=8'd68;
		data_a[19749]<=8'd51;
		data_a[19750]<=8'd49;
		data_a[19751]<=8'd55;
		data_a[19752]<=8'd36;
		data_a[19753]<=8'd44;
		data_a[19754]<=8'd58;
		data_a[19755]<=8'd47;
		data_a[19756]<=8'd37;
		data_a[19757]<=8'd46;
		data_a[19758]<=8'd46;
		data_a[19759]<=8'd37;
		data_a[19760]<=8'd41;
		data_a[19761]<=8'd36;
		data_a[19762]<=8'd42;
		data_a[19763]<=8'd39;
		data_a[19764]<=8'd41;
		data_a[19765]<=8'd41;
		data_a[19766]<=8'd45;
		data_a[19767]<=8'd36;
		data_a[19768]<=8'd39;
		data_a[19769]<=8'd45;
		data_a[19770]<=8'd43;
		data_a[19771]<=8'd39;
		data_a[19772]<=8'd43;
		data_a[19773]<=8'd40;
		data_a[19774]<=8'd47;
		data_a[19775]<=8'd54;
		data_a[19776]<=8'd97;
		data_a[19777]<=8'd112;
		data_a[19778]<=8'd128;
		data_a[19779]<=8'd127;
		data_a[19780]<=8'd132;
		data_a[19781]<=8'd134;
		data_a[19782]<=8'd124;
		data_a[19783]<=8'd114;
		data_a[19784]<=8'd100;
		data_a[19785]<=8'd71;
		data_a[19786]<=8'd74;
		data_a[19787]<=8'd77;
		data_a[19788]<=8'd80;
		data_a[19789]<=8'd89;
		data_a[19790]<=8'd92;
		data_a[19791]<=8'd114;
		data_a[19792]<=8'd120;
		data_a[19793]<=8'd112;
		data_a[19794]<=8'd103;
		data_a[19795]<=8'd97;
		data_a[19796]<=8'd94;
		data_a[19797]<=8'd100;
		data_a[19798]<=8'd95;
		data_a[19799]<=8'd89;
		data_a[19800]<=8'd254;
		data_a[19801]<=8'd91;
		data_a[19802]<=8'd92;
		data_a[19803]<=8'd86;
		data_a[19804]<=8'd81;
		data_a[19805]<=8'd66;
		data_a[19806]<=8'd58;
		data_a[19807]<=8'd52;
		data_a[19808]<=8'd49;
		data_a[19809]<=8'd65;
		data_a[19810]<=8'd78;
		data_a[19811]<=8'd80;
		data_a[19812]<=8'd75;
		data_a[19813]<=8'd70;
		data_a[19814]<=8'd98;
		data_a[19815]<=8'd104;
		data_a[19816]<=8'd97;
		data_a[19817]<=8'd86;
		data_a[19818]<=8'd75;
		data_a[19819]<=8'd108;
		data_a[19820]<=8'd173;
		data_a[19821]<=8'd177;
		data_a[19822]<=8'd171;
		data_a[19823]<=8'd168;
		data_a[19824]<=8'd191;
		data_a[19825]<=8'd175;
		data_a[19826]<=8'd180;
		data_a[19827]<=8'd185;
		data_a[19828]<=8'd194;
		data_a[19829]<=8'd193;
		data_a[19830]<=8'd200;
		data_a[19831]<=8'd184;
		data_a[19832]<=8'd133;
		data_a[19833]<=8'd129;
		data_a[19834]<=8'd108;
		data_a[19835]<=8'd65;
		data_a[19836]<=8'd63;
		data_a[19837]<=8'd55;
		data_a[19838]<=8'd63;
		data_a[19839]<=8'd81;
		data_a[19840]<=8'd85;
		data_a[19841]<=8'd84;
		data_a[19842]<=8'd86;
		data_a[19843]<=8'd96;
		data_a[19844]<=8'd94;
		data_a[19845]<=8'd101;
		data_a[19846]<=8'd107;
		data_a[19847]<=8'd99;
		data_a[19848]<=8'd96;
		data_a[19849]<=8'd93;
		data_a[19850]<=8'd83;
		data_a[19851]<=8'd71;
		data_a[19852]<=8'd68;
		data_a[19853]<=8'd70;
		data_a[19854]<=8'd62;
		data_a[19855]<=8'd99;
		data_a[19856]<=8'd122;
		data_a[19857]<=8'd138;
		data_a[19858]<=8'd235;
		data_a[19859]<=8'd232;
		data_a[19860]<=8'd232;
		data_a[19861]<=8'd236;
		data_a[19862]<=8'd235;
		data_a[19863]<=8'd238;
		data_a[19864]<=8'd235;
		data_a[19865]<=8'd234;
		data_a[19866]<=8'd235;
		data_a[19867]<=8'd236;
		data_a[19868]<=8'd235;
		data_a[19869]<=8'd234;
		data_a[19870]<=8'd234;
		data_a[19871]<=8'd235;
		data_a[19872]<=8'd236;
		data_a[19873]<=8'd234;
		data_a[19874]<=8'd234;
		data_a[19875]<=8'd235;
		data_a[19876]<=8'd235;
		data_a[19877]<=8'd239;
		data_a[19878]<=8'd242;
		data_a[19879]<=8'd241;
		data_a[19880]<=8'd241;
		data_a[19881]<=8'd241;
		data_a[19882]<=8'd242;
		data_a[19883]<=8'd242;
		data_a[19884]<=8'd241;
		data_a[19885]<=8'd241;
		data_a[19886]<=8'd241;
		data_a[19887]<=8'd241;
		data_a[19888]<=8'd237;
		data_a[19889]<=8'd241;
		data_a[19890]<=8'd243;
		data_a[19891]<=8'd235;
		data_a[19892]<=8'd228;
		data_a[19893]<=8'd247;
		data_a[19894]<=8'd195;
		data_a[19895]<=8'd54;
		data_a[19896]<=8'd93;
		data_a[19897]<=8'd59;
		data_a[19898]<=8'd58;
		data_a[19899]<=8'd49;
		data_a[19900]<=8'd48;
		data_a[19901]<=8'd49;
		data_a[19902]<=8'd49;
		data_a[19903]<=8'd40;
		data_a[19904]<=8'd47;
		data_a[19905]<=8'd44;
		data_a[19906]<=8'd51;
		data_a[19907]<=8'd42;
		data_a[19908]<=8'd35;
		data_a[19909]<=8'd41;
		data_a[19910]<=8'd38;
		data_a[19911]<=8'd39;
		data_a[19912]<=8'd38;
		data_a[19913]<=8'd39;
		data_a[19914]<=8'd43;
		data_a[19915]<=8'd41;
		data_a[19916]<=8'd44;
		data_a[19917]<=8'd39;
		data_a[19918]<=8'd41;
		data_a[19919]<=8'd44;
		data_a[19920]<=8'd42;
		data_a[19921]<=8'd41;
		data_a[19922]<=8'd39;
		data_a[19923]<=8'd46;
		data_a[19924]<=8'd46;
		data_a[19925]<=8'd83;
		data_a[19926]<=8'd104;
		data_a[19927]<=8'd114;
		data_a[19928]<=8'd128;
		data_a[19929]<=8'd129;
		data_a[19930]<=8'd133;
		data_a[19931]<=8'd132;
		data_a[19932]<=8'd121;
		data_a[19933]<=8'd115;
		data_a[19934]<=8'd100;
		data_a[19935]<=8'd70;
		data_a[19936]<=8'd71;
		data_a[19937]<=8'd73;
		data_a[19938]<=8'd81;
		data_a[19939]<=8'd81;
		data_a[19940]<=8'd97;
		data_a[19941]<=8'd110;
		data_a[19942]<=8'd121;
		data_a[19943]<=8'd118;
		data_a[19944]<=8'd103;
		data_a[19945]<=8'd95;
		data_a[19946]<=8'd93;
		data_a[19947]<=8'd96;
		data_a[19948]<=8'd94;
		data_a[19949]<=8'd90;
		data_a[19950]<=8'd255;
		data_a[19951]<=8'd84;
		data_a[19952]<=8'd87;
		data_a[19953]<=8'd91;
		data_a[19954]<=8'd88;
		data_a[19955]<=8'd67;
		data_a[19956]<=8'd60;
		data_a[19957]<=8'd54;
		data_a[19958]<=8'd47;
		data_a[19959]<=8'd75;
		data_a[19960]<=8'd73;
		data_a[19961]<=8'd76;
		data_a[19962]<=8'd77;
		data_a[19963]<=8'd144;
		data_a[19964]<=8'd248;
		data_a[19965]<=8'd230;
		data_a[19966]<=8'd66;
		data_a[19967]<=8'd79;
		data_a[19968]<=8'd80;
		data_a[19969]<=8'd90;
		data_a[19970]<=8'd153;
		data_a[19971]<=8'd165;
		data_a[19972]<=8'd174;
		data_a[19973]<=8'd180;
		data_a[19974]<=8'd179;
		data_a[19975]<=8'd149;
		data_a[19976]<=8'd185;
		data_a[19977]<=8'd186;
		data_a[19978]<=8'd197;
		data_a[19979]<=8'd194;
		data_a[19980]<=8'd197;
		data_a[19981]<=8'd176;
		data_a[19982]<=8'd134;
		data_a[19983]<=8'd127;
		data_a[19984]<=8'd109;
		data_a[19985]<=8'd73;
		data_a[19986]<=8'd66;
		data_a[19987]<=8'd60;
		data_a[19988]<=8'd60;
		data_a[19989]<=8'd71;
		data_a[19990]<=8'd77;
		data_a[19991]<=8'd78;
		data_a[19992]<=8'd74;
		data_a[19993]<=8'd90;
		data_a[19994]<=8'd92;
		data_a[19995]<=8'd98;
		data_a[19996]<=8'd103;
		data_a[19997]<=8'd90;
		data_a[19998]<=8'd82;
		data_a[19999]<=8'd81;
		data_a[20000]<=8'd79;
		data_a[20001]<=8'd66;
		data_a[20002]<=8'd68;
		data_a[20003]<=8'd63;
		data_a[20004]<=8'd71;
		data_a[20005]<=8'd106;
		data_a[20006]<=8'd115;
		data_a[20007]<=8'd146;
		data_a[20008]<=8'd235;
		data_a[20009]<=8'd233;
		data_a[20010]<=8'd237;
		data_a[20011]<=8'd236;
		data_a[20012]<=8'd234;
		data_a[20013]<=8'd234;
		data_a[20014]<=8'd234;
		data_a[20015]<=8'd234;
		data_a[20016]<=8'd235;
		data_a[20017]<=8'd236;
		data_a[20018]<=8'd235;
		data_a[20019]<=8'd234;
		data_a[20020]<=8'd234;
		data_a[20021]<=8'd235;
		data_a[20022]<=8'd234;
		data_a[20023]<=8'd234;
		data_a[20024]<=8'd233;
		data_a[20025]<=8'd236;
		data_a[20026]<=8'd235;
		data_a[20027]<=8'd240;
		data_a[20028]<=8'd241;
		data_a[20029]<=8'd239;
		data_a[20030]<=8'd241;
		data_a[20031]<=8'd241;
		data_a[20032]<=8'd242;
		data_a[20033]<=8'd242;
		data_a[20034]<=8'd242;
		data_a[20035]<=8'd240;
		data_a[20036]<=8'd240;
		data_a[20037]<=8'd240;
		data_a[20038]<=8'd245;
		data_a[20039]<=8'd236;
		data_a[20040]<=8'd241;
		data_a[20041]<=8'd242;
		data_a[20042]<=8'd246;
		data_a[20043]<=8'd248;
		data_a[20044]<=8'd241;
		data_a[20045]<=8'd110;
		data_a[20046]<=8'd162;
		data_a[20047]<=8'd43;
		data_a[20048]<=8'd47;
		data_a[20049]<=8'd56;
		data_a[20050]<=8'd50;
		data_a[20051]<=8'd52;
		data_a[20052]<=8'd43;
		data_a[20053]<=8'd41;
		data_a[20054]<=8'd41;
		data_a[20055]<=8'd46;
		data_a[20056]<=8'd39;
		data_a[20057]<=8'd36;
		data_a[20058]<=8'd37;
		data_a[20059]<=8'd41;
		data_a[20060]<=8'd44;
		data_a[20061]<=8'd30;
		data_a[20062]<=8'd40;
		data_a[20063]<=8'd41;
		data_a[20064]<=8'd42;
		data_a[20065]<=8'd41;
		data_a[20066]<=8'd42;
		data_a[20067]<=8'd38;
		data_a[20068]<=8'd40;
		data_a[20069]<=8'd44;
		data_a[20070]<=8'd47;
		data_a[20071]<=8'd43;
		data_a[20072]<=8'd44;
		data_a[20073]<=8'd39;
		data_a[20074]<=8'd64;
		data_a[20075]<=8'd98;
		data_a[20076]<=8'd108;
		data_a[20077]<=8'd116;
		data_a[20078]<=8'd127;
		data_a[20079]<=8'd128;
		data_a[20080]<=8'd131;
		data_a[20081]<=8'd130;
		data_a[20082]<=8'd119;
		data_a[20083]<=8'd116;
		data_a[20084]<=8'd97;
		data_a[20085]<=8'd69;
		data_a[20086]<=8'd72;
		data_a[20087]<=8'd76;
		data_a[20088]<=8'd79;
		data_a[20089]<=8'd81;
		data_a[20090]<=8'd95;
		data_a[20091]<=8'd108;
		data_a[20092]<=8'd115;
		data_a[20093]<=8'd122;
		data_a[20094]<=8'd102;
		data_a[20095]<=8'd94;
		data_a[20096]<=8'd92;
		data_a[20097]<=8'd92;
		data_a[20098]<=8'd94;
		data_a[20099]<=8'd91;
		data_a[20100]<=8'd255;
		data_a[20101]<=8'd90;
		data_a[20102]<=8'd90;
		data_a[20103]<=8'd86;
		data_a[20104]<=8'd80;
		data_a[20105]<=8'd62;
		data_a[20106]<=8'd60;
		data_a[20107]<=8'd58;
		data_a[20108]<=8'd51;
		data_a[20109]<=8'd70;
		data_a[20110]<=8'd77;
		data_a[20111]<=8'd81;
		data_a[20112]<=8'd178;
		data_a[20113]<=8'd243;
		data_a[20114]<=8'd245;
		data_a[20115]<=8'd245;
		data_a[20116]<=8'd227;
		data_a[20117]<=8'd57;
		data_a[20118]<=8'd64;
		data_a[20119]<=8'd76;
		data_a[20120]<=8'd146;
		data_a[20121]<=8'd149;
		data_a[20122]<=8'd130;
		data_a[20123]<=8'd115;
		data_a[20124]<=8'd134;
		data_a[20125]<=8'd116;
		data_a[20126]<=8'd190;
		data_a[20127]<=8'd187;
		data_a[20128]<=8'd189;
		data_a[20129]<=8'd198;
		data_a[20130]<=8'd200;
		data_a[20131]<=8'd153;
		data_a[20132]<=8'd136;
		data_a[20133]<=8'd132;
		data_a[20134]<=8'd122;
		data_a[20135]<=8'd92;
		data_a[20136]<=8'd68;
		data_a[20137]<=8'd53;
		data_a[20138]<=8'd56;
		data_a[20139]<=8'd63;
		data_a[20140]<=8'd69;
		data_a[20141]<=8'd70;
		data_a[20142]<=8'd69;
		data_a[20143]<=8'd80;
		data_a[20144]<=8'd88;
		data_a[20145]<=8'd91;
		data_a[20146]<=8'd90;
		data_a[20147]<=8'd79;
		data_a[20148]<=8'd75;
		data_a[20149]<=8'd73;
		data_a[20150]<=8'd66;
		data_a[20151]<=8'd60;
		data_a[20152]<=8'd59;
		data_a[20153]<=8'd62;
		data_a[20154]<=8'd94;
		data_a[20155]<=8'd110;
		data_a[20156]<=8'd122;
		data_a[20157]<=8'd167;
		data_a[20158]<=8'd237;
		data_a[20159]<=8'd232;
		data_a[20160]<=8'd234;
		data_a[20161]<=8'd234;
		data_a[20162]<=8'd233;
		data_a[20163]<=8'd234;
		data_a[20164]<=8'd234;
		data_a[20165]<=8'd234;
		data_a[20166]<=8'd235;
		data_a[20167]<=8'd235;
		data_a[20168]<=8'd235;
		data_a[20169]<=8'd234;
		data_a[20170]<=8'd234;
		data_a[20171]<=8'd235;
		data_a[20172]<=8'd234;
		data_a[20173]<=8'd234;
		data_a[20174]<=8'd233;
		data_a[20175]<=8'd237;
		data_a[20176]<=8'd235;
		data_a[20177]<=8'd241;
		data_a[20178]<=8'd240;
		data_a[20179]<=8'd238;
		data_a[20180]<=8'd241;
		data_a[20181]<=8'd240;
		data_a[20182]<=8'd241;
		data_a[20183]<=8'd242;
		data_a[20184]<=8'd241;
		data_a[20185]<=8'd240;
		data_a[20186]<=8'd240;
		data_a[20187]<=8'd242;
		data_a[20188]<=8'd242;
		data_a[20189]<=8'd241;
		data_a[20190]<=8'd239;
		data_a[20191]<=8'd238;
		data_a[20192]<=8'd235;
		data_a[20193]<=8'd242;
		data_a[20194]<=8'd250;
		data_a[20195]<=8'd170;
		data_a[20196]<=8'd89;
		data_a[20197]<=8'd67;
		data_a[20198]<=8'd49;
		data_a[20199]<=8'd42;
		data_a[20200]<=8'd45;
		data_a[20201]<=8'd44;
		data_a[20202]<=8'd45;
		data_a[20203]<=8'd42;
		data_a[20204]<=8'd42;
		data_a[20205]<=8'd35;
		data_a[20206]<=8'd38;
		data_a[20207]<=8'd41;
		data_a[20208]<=8'd39;
		data_a[20209]<=8'd34;
		data_a[20210]<=8'd32;
		data_a[20211]<=8'd45;
		data_a[20212]<=8'd40;
		data_a[20213]<=8'd44;
		data_a[20214]<=8'd42;
		data_a[20215]<=8'd40;
		data_a[20216]<=8'd39;
		data_a[20217]<=8'd41;
		data_a[20218]<=8'd41;
		data_a[20219]<=8'd43;
		data_a[20220]<=8'd43;
		data_a[20221]<=8'd51;
		data_a[20222]<=8'd61;
		data_a[20223]<=8'd67;
		data_a[20224]<=8'd80;
		data_a[20225]<=8'd104;
		data_a[20226]<=8'd104;
		data_a[20227]<=8'd120;
		data_a[20228]<=8'd125;
		data_a[20229]<=8'd126;
		data_a[20230]<=8'd127;
		data_a[20231]<=8'd127;
		data_a[20232]<=8'd118;
		data_a[20233]<=8'd114;
		data_a[20234]<=8'd92;
		data_a[20235]<=8'd70;
		data_a[20236]<=8'd72;
		data_a[20237]<=8'd74;
		data_a[20238]<=8'd74;
		data_a[20239]<=8'd83;
		data_a[20240]<=8'd90;
		data_a[20241]<=8'd109;
		data_a[20242]<=8'd112;
		data_a[20243]<=8'd125;
		data_a[20244]<=8'd99;
		data_a[20245]<=8'd95;
		data_a[20246]<=8'd94;
		data_a[20247]<=8'd89;
		data_a[20248]<=8'd93;
		data_a[20249]<=8'd90;
		data_a[20250]<=8'd254;
		data_a[20251]<=8'd89;
		data_a[20252]<=8'd86;
		data_a[20253]<=8'd87;
		data_a[20254]<=8'd87;
		data_a[20255]<=8'd64;
		data_a[20256]<=8'd56;
		data_a[20257]<=8'd56;
		data_a[20258]<=8'd52;
		data_a[20259]<=8'd73;
		data_a[20260]<=8'd79;
		data_a[20261]<=8'd109;
		data_a[20262]<=8'd228;
		data_a[20263]<=8'd239;
		data_a[20264]<=8'd247;
		data_a[20265]<=8'd245;
		data_a[20266]<=8'd232;
		data_a[20267]<=8'd147;
		data_a[20268]<=8'd71;
		data_a[20269]<=8'd73;
		data_a[20270]<=8'd91;
		data_a[20271]<=8'd132;
		data_a[20272]<=8'd131;
		data_a[20273]<=8'd104;
		data_a[20274]<=8'd107;
		data_a[20275]<=8'd144;
		data_a[20276]<=8'd106;
		data_a[20277]<=8'd182;
		data_a[20278]<=8'd192;
		data_a[20279]<=8'd196;
		data_a[20280]<=8'd191;
		data_a[20281]<=8'd154;
		data_a[20282]<=8'd138;
		data_a[20283]<=8'd132;
		data_a[20284]<=8'd125;
		data_a[20285]<=8'd103;
		data_a[20286]<=8'd80;
		data_a[20287]<=8'd57;
		data_a[20288]<=8'd65;
		data_a[20289]<=8'd60;
		data_a[20290]<=8'd63;
		data_a[20291]<=8'd63;
		data_a[20292]<=8'd70;
		data_a[20293]<=8'd73;
		data_a[20294]<=8'd83;
		data_a[20295]<=8'd83;
		data_a[20296]<=8'd80;
		data_a[20297]<=8'd73;
		data_a[20298]<=8'd68;
		data_a[20299]<=8'd67;
		data_a[20300]<=8'd64;
		data_a[20301]<=8'd57;
		data_a[20302]<=8'd60;
		data_a[20303]<=8'd81;
		data_a[20304]<=8'd96;
		data_a[20305]<=8'd112;
		data_a[20306]<=8'd122;
		data_a[20307]<=8'd168;
		data_a[20308]<=8'd231;
		data_a[20309]<=8'd230;
		data_a[20310]<=8'd230;
		data_a[20311]<=8'd235;
		data_a[20312]<=8'd233;
		data_a[20313]<=8'd236;
		data_a[20314]<=8'd234;
		data_a[20315]<=8'd234;
		data_a[20316]<=8'd235;
		data_a[20317]<=8'd235;
		data_a[20318]<=8'd235;
		data_a[20319]<=8'd234;
		data_a[20320]<=8'd234;
		data_a[20321]<=8'd234;
		data_a[20322]<=8'd236;
		data_a[20323]<=8'd235;
		data_a[20324]<=8'd232;
		data_a[20325]<=8'd236;
		data_a[20326]<=8'd233;
		data_a[20327]<=8'd240;
		data_a[20328]<=8'd240;
		data_a[20329]<=8'd239;
		data_a[20330]<=8'd240;
		data_a[20331]<=8'd239;
		data_a[20332]<=8'd240;
		data_a[20333]<=8'd241;
		data_a[20334]<=8'd241;
		data_a[20335]<=8'd241;
		data_a[20336]<=8'd242;
		data_a[20337]<=8'd244;
		data_a[20338]<=8'd238;
		data_a[20339]<=8'd240;
		data_a[20340]<=8'd237;
		data_a[20341]<=8'd239;
		data_a[20342]<=8'd247;
		data_a[20343]<=8'd245;
		data_a[20344]<=8'd235;
		data_a[20345]<=8'd238;
		data_a[20346]<=8'd132;
		data_a[20347]<=8'd68;
		data_a[20348]<=8'd49;
		data_a[20349]<=8'd53;
		data_a[20350]<=8'd46;
		data_a[20351]<=8'd52;
		data_a[20352]<=8'd41;
		data_a[20353]<=8'd36;
		data_a[20354]<=8'd37;
		data_a[20355]<=8'd41;
		data_a[20356]<=8'd37;
		data_a[20357]<=8'd34;
		data_a[20358]<=8'd37;
		data_a[20359]<=8'd38;
		data_a[20360]<=8'd39;
		data_a[20361]<=8'd41;
		data_a[20362]<=8'd40;
		data_a[20363]<=8'd42;
		data_a[20364]<=8'd39;
		data_a[20365]<=8'd43;
		data_a[20366]<=8'd41;
		data_a[20367]<=8'd43;
		data_a[20368]<=8'd42;
		data_a[20369]<=8'd48;
		data_a[20370]<=8'd58;
		data_a[20371]<=8'd55;
		data_a[20372]<=8'd75;
		data_a[20373]<=8'd83;
		data_a[20374]<=8'd96;
		data_a[20375]<=8'd104;
		data_a[20376]<=8'd113;
		data_a[20377]<=8'd121;
		data_a[20378]<=8'd125;
		data_a[20379]<=8'd124;
		data_a[20380]<=8'd123;
		data_a[20381]<=8'd125;
		data_a[20382]<=8'd118;
		data_a[20383]<=8'd112;
		data_a[20384]<=8'd88;
		data_a[20385]<=8'd70;
		data_a[20386]<=8'd77;
		data_a[20387]<=8'd70;
		data_a[20388]<=8'd77;
		data_a[20389]<=8'd80;
		data_a[20390]<=8'd92;
		data_a[20391]<=8'd103;
		data_a[20392]<=8'd113;
		data_a[20393]<=8'd122;
		data_a[20394]<=8'd97;
		data_a[20395]<=8'd96;
		data_a[20396]<=8'd95;
		data_a[20397]<=8'd87;
		data_a[20398]<=8'd92;
		data_a[20399]<=8'd88;
		data_a[20400]<=8'd254;
		data_a[20401]<=8'd90;
		data_a[20402]<=8'd88;
		data_a[20403]<=8'd86;
		data_a[20404]<=8'd86;
		data_a[20405]<=8'd64;
		data_a[20406]<=8'd61;
		data_a[20407]<=8'd56;
		data_a[20408]<=8'd49;
		data_a[20409]<=8'd72;
		data_a[20410]<=8'd77;
		data_a[20411]<=8'd250;
		data_a[20412]<=8'd209;
		data_a[20413]<=8'd230;
		data_a[20414]<=8'd228;
		data_a[20415]<=8'd225;
		data_a[20416]<=8'd208;
		data_a[20417]<=8'd53;
		data_a[20418]<=8'd65;
		data_a[20419]<=8'd65;
		data_a[20420]<=8'd76;
		data_a[20421]<=8'd132;
		data_a[20422]<=8'd120;
		data_a[20423]<=8'd108;
		data_a[20424]<=8'd92;
		data_a[20425]<=8'd100;
		data_a[20426]<=8'd133;
		data_a[20427]<=8'd72;
		data_a[20428]<=8'd196;
		data_a[20429]<=8'd213;
		data_a[20430]<=8'd151;
		data_a[20431]<=8'd157;
		data_a[20432]<=8'd140;
		data_a[20433]<=8'd131;
		data_a[20434]<=8'd128;
		data_a[20435]<=8'd115;
		data_a[20436]<=8'd97;
		data_a[20437]<=8'd71;
		data_a[20438]<=8'd61;
		data_a[20439]<=8'd57;
		data_a[20440]<=8'd62;
		data_a[20441]<=8'd64;
		data_a[20442]<=8'd65;
		data_a[20443]<=8'd66;
		data_a[20444]<=8'd75;
		data_a[20445]<=8'd75;
		data_a[20446]<=8'd76;
		data_a[20447]<=8'd67;
		data_a[20448]<=8'd65;
		data_a[20449]<=8'd61;
		data_a[20450]<=8'd55;
		data_a[20451]<=8'd55;
		data_a[20452]<=8'd67;
		data_a[20453]<=8'd86;
		data_a[20454]<=8'd102;
		data_a[20455]<=8'd108;
		data_a[20456]<=8'd122;
		data_a[20457]<=8'd172;
		data_a[20458]<=8'd235;
		data_a[20459]<=8'd231;
		data_a[20460]<=8'd231;
		data_a[20461]<=8'd237;
		data_a[20462]<=8'd228;
		data_a[20463]<=8'd237;
		data_a[20464]<=8'd237;
		data_a[20465]<=8'd234;
		data_a[20466]<=8'd237;
		data_a[20467]<=8'd234;
		data_a[20468]<=8'd234;
		data_a[20469]<=8'd238;
		data_a[20470]<=8'd236;
		data_a[20471]<=8'd236;
		data_a[20472]<=8'd237;
		data_a[20473]<=8'd235;
		data_a[20474]<=8'd235;
		data_a[20475]<=8'd235;
		data_a[20476]<=8'd233;
		data_a[20477]<=8'd235;
		data_a[20478]<=8'd238;
		data_a[20479]<=8'd238;
		data_a[20480]<=8'd242;
		data_a[20481]<=8'd239;
		data_a[20482]<=8'd240;
		data_a[20483]<=8'd240;
		data_a[20484]<=8'd240;
		data_a[20485]<=8'd241;
		data_a[20486]<=8'd241;
		data_a[20487]<=8'd239;
		data_a[20488]<=8'd242;
		data_a[20489]<=8'd238;
		data_a[20490]<=8'd239;
		data_a[20491]<=8'd239;
		data_a[20492]<=8'd243;
		data_a[20493]<=8'd241;
		data_a[20494]<=8'd239;
		data_a[20495]<=8'd232;
		data_a[20496]<=8'd183;
		data_a[20497]<=8'd61;
		data_a[20498]<=8'd52;
		data_a[20499]<=8'd46;
		data_a[20500]<=8'd42;
		data_a[20501]<=8'd52;
		data_a[20502]<=8'd45;
		data_a[20503]<=8'd39;
		data_a[20504]<=8'd40;
		data_a[20505]<=8'd41;
		data_a[20506]<=8'd34;
		data_a[20507]<=8'd35;
		data_a[20508]<=8'd36;
		data_a[20509]<=8'd36;
		data_a[20510]<=8'd44;
		data_a[20511]<=8'd43;
		data_a[20512]<=8'd37;
		data_a[20513]<=8'd41;
		data_a[20514]<=8'd39;
		data_a[20515]<=8'd42;
		data_a[20516]<=8'd45;
		data_a[20517]<=8'd36;
		data_a[20518]<=8'd51;
		data_a[20519]<=8'd62;
		data_a[20520]<=8'd68;
		data_a[20521]<=8'd80;
		data_a[20522]<=8'd86;
		data_a[20523]<=8'd92;
		data_a[20524]<=8'd102;
		data_a[20525]<=8'd108;
		data_a[20526]<=8'd112;
		data_a[20527]<=8'd122;
		data_a[20528]<=8'd124;
		data_a[20529]<=8'd121;
		data_a[20530]<=8'd125;
		data_a[20531]<=8'd120;
		data_a[20532]<=8'd114;
		data_a[20533]<=8'd109;
		data_a[20534]<=8'd89;
		data_a[20535]<=8'd69;
		data_a[20536]<=8'd72;
		data_a[20537]<=8'd74;
		data_a[20538]<=8'd71;
		data_a[20539]<=8'd78;
		data_a[20540]<=8'd90;
		data_a[20541]<=8'd98;
		data_a[20542]<=8'd114;
		data_a[20543]<=8'd120;
		data_a[20544]<=8'd96;
		data_a[20545]<=8'd93;
		data_a[20546]<=8'd97;
		data_a[20547]<=8'd88;
		data_a[20548]<=8'd91;
		data_a[20549]<=8'd90;
		data_a[20550]<=8'd253;
		data_a[20551]<=8'd87;
		data_a[20552]<=8'd93;
		data_a[20553]<=8'd83;
		data_a[20554]<=8'd84;
		data_a[20555]<=8'd71;
		data_a[20556]<=8'd50;
		data_a[20557]<=8'd68;
		data_a[20558]<=8'd53;
		data_a[20559]<=8'd66;
		data_a[20560]<=8'd161;
		data_a[20561]<=8'd214;
		data_a[20562]<=8'd214;
		data_a[20563]<=8'd234;
		data_a[20564]<=8'd232;
		data_a[20565]<=8'd172;
		data_a[20566]<=8'd39;
		data_a[20567]<=8'd62;
		data_a[20568]<=8'd60;
		data_a[20569]<=8'd67;
		data_a[20570]<=8'd72;
		data_a[20571]<=8'd101;
		data_a[20572]<=8'd100;
		data_a[20573]<=8'd97;
		data_a[20574]<=8'd69;
		data_a[20575]<=8'd80;
		data_a[20576]<=8'd86;
		data_a[20577]<=8'd114;
		data_a[20578]<=8'd229;
		data_a[20579]<=8'd183;
		data_a[20580]<=8'd151;
		data_a[20581]<=8'd151;
		data_a[20582]<=8'd141;
		data_a[20583]<=8'd131;
		data_a[20584]<=8'd126;
		data_a[20585]<=8'd119;
		data_a[20586]<=8'd113;
		data_a[20587]<=8'd95;
		data_a[20588]<=8'd79;
		data_a[20589]<=8'd63;
		data_a[20590]<=8'd57;
		data_a[20591]<=8'd57;
		data_a[20592]<=8'd63;
		data_a[20593]<=8'd67;
		data_a[20594]<=8'd70;
		data_a[20595]<=8'd72;
		data_a[20596]<=8'd65;
		data_a[20597]<=8'd63;
		data_a[20598]<=8'd63;
		data_a[20599]<=8'd56;
		data_a[20600]<=8'd53;
		data_a[20601]<=8'd63;
		data_a[20602]<=8'd81;
		data_a[20603]<=8'd97;
		data_a[20604]<=8'd107;
		data_a[20605]<=8'd111;
		data_a[20606]<=8'd123;
		data_a[20607]<=8'd167;
		data_a[20608]<=8'd233;
		data_a[20609]<=8'd231;
		data_a[20610]<=8'd228;
		data_a[20611]<=8'd236;
		data_a[20612]<=8'd238;
		data_a[20613]<=8'd230;
		data_a[20614]<=8'd229;
		data_a[20615]<=8'd235;
		data_a[20616]<=8'd235;
		data_a[20617]<=8'd232;
		data_a[20618]<=8'd238;
		data_a[20619]<=8'd231;
		data_a[20620]<=8'd229;
		data_a[20621]<=8'd240;
		data_a[20622]<=8'd236;
		data_a[20623]<=8'd234;
		data_a[20624]<=8'd234;
		data_a[20625]<=8'd234;
		data_a[20626]<=8'd234;
		data_a[20627]<=8'd236;
		data_a[20628]<=8'd239;
		data_a[20629]<=8'd239;
		data_a[20630]<=8'd241;
		data_a[20631]<=8'd239;
		data_a[20632]<=8'd239;
		data_a[20633]<=8'd240;
		data_a[20634]<=8'd239;
		data_a[20635]<=8'd240;
		data_a[20636]<=8'd241;
		data_a[20637]<=8'd239;
		data_a[20638]<=8'd241;
		data_a[20639]<=8'd238;
		data_a[20640]<=8'd239;
		data_a[20641]<=8'd238;
		data_a[20642]<=8'd243;
		data_a[20643]<=8'd242;
		data_a[20644]<=8'd241;
		data_a[20645]<=8'd236;
		data_a[20646]<=8'd249;
		data_a[20647]<=8'd58;
		data_a[20648]<=8'd46;
		data_a[20649]<=8'd47;
		data_a[20650]<=8'd46;
		data_a[20651]<=8'd47;
		data_a[20652]<=8'd40;
		data_a[20653]<=8'd44;
		data_a[20654]<=8'd41;
		data_a[20655]<=8'd36;
		data_a[20656]<=8'd39;
		data_a[20657]<=8'd38;
		data_a[20658]<=8'd39;
		data_a[20659]<=8'd43;
		data_a[20660]<=8'd37;
		data_a[20661]<=8'd38;
		data_a[20662]<=8'd39;
		data_a[20663]<=8'd38;
		data_a[20664]<=8'd38;
		data_a[20665]<=8'd45;
		data_a[20666]<=8'd43;
		data_a[20667]<=8'd58;
		data_a[20668]<=8'd72;
		data_a[20669]<=8'd73;
		data_a[20670]<=8'd76;
		data_a[20671]<=8'd82;
		data_a[20672]<=8'd90;
		data_a[20673]<=8'd98;
		data_a[20674]<=8'd105;
		data_a[20675]<=8'd110;
		data_a[20676]<=8'd117;
		data_a[20677]<=8'd123;
		data_a[20678]<=8'd125;
		data_a[20679]<=8'd123;
		data_a[20680]<=8'd125;
		data_a[20681]<=8'd120;
		data_a[20682]<=8'd114;
		data_a[20683]<=8'd109;
		data_a[20684]<=8'd87;
		data_a[20685]<=8'd66;
		data_a[20686]<=8'd68;
		data_a[20687]<=8'd63;
		data_a[20688]<=8'd75;
		data_a[20689]<=8'd81;
		data_a[20690]<=8'd89;
		data_a[20691]<=8'd101;
		data_a[20692]<=8'd107;
		data_a[20693]<=8'd117;
		data_a[20694]<=8'd103;
		data_a[20695]<=8'd93;
		data_a[20696]<=8'd95;
		data_a[20697]<=8'd90;
		data_a[20698]<=8'd88;
		data_a[20699]<=8'd86;
		data_a[20700]<=8'd254;
		data_a[20701]<=8'd93;
		data_a[20702]<=8'd79;
		data_a[20703]<=8'd88;
		data_a[20704]<=8'd83;
		data_a[20705]<=8'd58;
		data_a[20706]<=8'd53;
		data_a[20707]<=8'd71;
		data_a[20708]<=8'd51;
		data_a[20709]<=8'd79;
		data_a[20710]<=8'd244;
		data_a[20711]<=8'd182;
		data_a[20712]<=8'd209;
		data_a[20713]<=8'd216;
		data_a[20714]<=8'd179;
		data_a[20715]<=8'd45;
		data_a[20716]<=8'd60;
		data_a[20717]<=8'd61;
		data_a[20718]<=8'd66;
		data_a[20719]<=8'd66;
		data_a[20720]<=8'd65;
		data_a[20721]<=8'd86;
		data_a[20722]<=8'd90;
		data_a[20723]<=8'd64;
		data_a[20724]<=8'd60;
		data_a[20725]<=8'd113;
		data_a[20726]<=8'd200;
		data_a[20727]<=8'd218;
		data_a[20728]<=8'd214;
		data_a[20729]<=8'd66;
		data_a[20730]<=8'd174;
		data_a[20731]<=8'd158;
		data_a[20732]<=8'd141;
		data_a[20733]<=8'd134;
		data_a[20734]<=8'd129;
		data_a[20735]<=8'd122;
		data_a[20736]<=8'd119;
		data_a[20737]<=8'd111;
		data_a[20738]<=8'd99;
		data_a[20739]<=8'd84;
		data_a[20740]<=8'd77;
		data_a[20741]<=8'd61;
		data_a[20742]<=8'd56;
		data_a[20743]<=8'd56;
		data_a[20744]<=8'd57;
		data_a[20745]<=8'd64;
		data_a[20746]<=8'd53;
		data_a[20747]<=8'd58;
		data_a[20748]<=8'd54;
		data_a[20749]<=8'd54;
		data_a[20750]<=8'd63;
		data_a[20751]<=8'd78;
		data_a[20752]<=8'd90;
		data_a[20753]<=8'd95;
		data_a[20754]<=8'd102;
		data_a[20755]<=8'd110;
		data_a[20756]<=8'd125;
		data_a[20757]<=8'd149;
		data_a[20758]<=8'd232;
		data_a[20759]<=8'd238;
		data_a[20760]<=8'd219;
		data_a[20761]<=8'd174;
		data_a[20762]<=8'd174;
		data_a[20763]<=8'd234;
		data_a[20764]<=8'd238;
		data_a[20765]<=8'd232;
		data_a[20766]<=8'd238;
		data_a[20767]<=8'd236;
		data_a[20768]<=8'd234;
		data_a[20769]<=8'd241;
		data_a[20770]<=8'd232;
		data_a[20771]<=8'd237;
		data_a[20772]<=8'd236;
		data_a[20773]<=8'd233;
		data_a[20774]<=8'd233;
		data_a[20775]<=8'd234;
		data_a[20776]<=8'd234;
		data_a[20777]<=8'd236;
		data_a[20778]<=8'd239;
		data_a[20779]<=8'd238;
		data_a[20780]<=8'd240;
		data_a[20781]<=8'd238;
		data_a[20782]<=8'd238;
		data_a[20783]<=8'd239;
		data_a[20784]<=8'd239;
		data_a[20785]<=8'd240;
		data_a[20786]<=8'd241;
		data_a[20787]<=8'd239;
		data_a[20788]<=8'd240;
		data_a[20789]<=8'd236;
		data_a[20790]<=8'd237;
		data_a[20791]<=8'd237;
		data_a[20792]<=8'd243;
		data_a[20793]<=8'd242;
		data_a[20794]<=8'd242;
		data_a[20795]<=8'd239;
		data_a[20796]<=8'd192;
		data_a[20797]<=8'd164;
		data_a[20798]<=8'd50;
		data_a[20799]<=8'd49;
		data_a[20800]<=8'd47;
		data_a[20801]<=8'd47;
		data_a[20802]<=8'd50;
		data_a[20803]<=8'd36;
		data_a[20804]<=8'd41;
		data_a[20805]<=8'd42;
		data_a[20806]<=8'd48;
		data_a[20807]<=8'd43;
		data_a[20808]<=8'd39;
		data_a[20809]<=8'd40;
		data_a[20810]<=8'd41;
		data_a[20811]<=8'd48;
		data_a[20812]<=8'd39;
		data_a[20813]<=8'd41;
		data_a[20814]<=8'd41;
		data_a[20815]<=8'd48;
		data_a[20816]<=8'd60;
		data_a[20817]<=8'd80;
		data_a[20818]<=8'd82;
		data_a[20819]<=8'd84;
		data_a[20820]<=8'd87;
		data_a[20821]<=8'd88;
		data_a[20822]<=8'd96;
		data_a[20823]<=8'd103;
		data_a[20824]<=8'd106;
		data_a[20825]<=8'd113;
		data_a[20826]<=8'd121;
		data_a[20827]<=8'd123;
		data_a[20828]<=8'd124;
		data_a[20829]<=8'd124;
		data_a[20830]<=8'd124;
		data_a[20831]<=8'd118;
		data_a[20832]<=8'd113;
		data_a[20833]<=8'd107;
		data_a[20834]<=8'd86;
		data_a[20835]<=8'd63;
		data_a[20836]<=8'd71;
		data_a[20837]<=8'd67;
		data_a[20838]<=8'd70;
		data_a[20839]<=8'd81;
		data_a[20840]<=8'd85;
		data_a[20841]<=8'd89;
		data_a[20842]<=8'd97;
		data_a[20843]<=8'd101;
		data_a[20844]<=8'd111;
		data_a[20845]<=8'd95;
		data_a[20846]<=8'd95;
		data_a[20847]<=8'd93;
		data_a[20848]<=8'd88;
		data_a[20849]<=8'd85;
		data_a[20850]<=8'd254;
		data_a[20851]<=8'd87;
		data_a[20852]<=8'd87;
		data_a[20853]<=8'd90;
		data_a[20854]<=8'd79;
		data_a[20855]<=8'd69;
		data_a[20856]<=8'd63;
		data_a[20857]<=8'd68;
		data_a[20858]<=8'd52;
		data_a[20859]<=8'd107;
		data_a[20860]<=8'd210;
		data_a[20861]<=8'd162;
		data_a[20862]<=8'd204;
		data_a[20863]<=8'd198;
		data_a[20864]<=8'd70;
		data_a[20865]<=8'd78;
		data_a[20866]<=8'd75;
		data_a[20867]<=8'd68;
		data_a[20868]<=8'd68;
		data_a[20869]<=8'd58;
		data_a[20870]<=8'd62;
		data_a[20871]<=8'd65;
		data_a[20872]<=8'd58;
		data_a[20873]<=8'd39;
		data_a[20874]<=8'd106;
		data_a[20875]<=8'd208;
		data_a[20876]<=8'd209;
		data_a[20877]<=8'd207;
		data_a[20878]<=8'd202;
		data_a[20879]<=8'd110;
		data_a[20880]<=8'd161;
		data_a[20881]<=8'd149;
		data_a[20882]<=8'd141;
		data_a[20883]<=8'd137;
		data_a[20884]<=8'd132;
		data_a[20885]<=8'd123;
		data_a[20886]<=8'd117;
		data_a[20887]<=8'd114;
		data_a[20888]<=8'd110;
		data_a[20889]<=8'd101;
		data_a[20890]<=8'd100;
		data_a[20891]<=8'd90;
		data_a[20892]<=8'd87;
		data_a[20893]<=8'd82;
		data_a[20894]<=8'd74;
		data_a[20895]<=8'd73;
		data_a[20896]<=8'd68;
		data_a[20897]<=8'd77;
		data_a[20898]<=8'd65;
		data_a[20899]<=8'd70;
		data_a[20900]<=8'd81;
		data_a[20901]<=8'd93;
		data_a[20902]<=8'd95;
		data_a[20903]<=8'd93;
		data_a[20904]<=8'd100;
		data_a[20905]<=8'd111;
		data_a[20906]<=8'd120;
		data_a[20907]<=8'd151;
		data_a[20908]<=8'd171;
		data_a[20909]<=8'd150;
		data_a[20910]<=8'd122;
		data_a[20911]<=8'd103;
		data_a[20912]<=8'd166;
		data_a[20913]<=8'd170;
		data_a[20914]<=8'd234;
		data_a[20915]<=8'd234;
		data_a[20916]<=8'd231;
		data_a[20917]<=8'd230;
		data_a[20918]<=8'd235;
		data_a[20919]<=8'd230;
		data_a[20920]<=8'd235;
		data_a[20921]<=8'd239;
		data_a[20922]<=8'd236;
		data_a[20923]<=8'd233;
		data_a[20924]<=8'd233;
		data_a[20925]<=8'd233;
		data_a[20926]<=8'd233;
		data_a[20927]<=8'd235;
		data_a[20928]<=8'd238;
		data_a[20929]<=8'd237;
		data_a[20930]<=8'd239;
		data_a[20931]<=8'd237;
		data_a[20932]<=8'd238;
		data_a[20933]<=8'd239;
		data_a[20934]<=8'd239;
		data_a[20935]<=8'd240;
		data_a[20936]<=8'd241;
		data_a[20937]<=8'd239;
		data_a[20938]<=8'd240;
		data_a[20939]<=8'd236;
		data_a[20940]<=8'd236;
		data_a[20941]<=8'd236;
		data_a[20942]<=8'd244;
		data_a[20943]<=8'd243;
		data_a[20944]<=8'd242;
		data_a[20945]<=8'd240;
		data_a[20946]<=8'd249;
		data_a[20947]<=8'd236;
		data_a[20948]<=8'd52;
		data_a[20949]<=8'd48;
		data_a[20950]<=8'd49;
		data_a[20951]<=8'd41;
		data_a[20952]<=8'd38;
		data_a[20953]<=8'd45;
		data_a[20954]<=8'd36;
		data_a[20955]<=8'd39;
		data_a[20956]<=8'd36;
		data_a[20957]<=8'd40;
		data_a[20958]<=8'd44;
		data_a[20959]<=8'd48;
		data_a[20960]<=8'd59;
		data_a[20961]<=8'd61;
		data_a[20962]<=8'd56;
		data_a[20963]<=8'd53;
		data_a[20964]<=8'd60;
		data_a[20965]<=8'd62;
		data_a[20966]<=8'd81;
		data_a[20967]<=8'd87;
		data_a[20968]<=8'd84;
		data_a[20969]<=8'd90;
		data_a[20970]<=8'd94;
		data_a[20971]<=8'd97;
		data_a[20972]<=8'd101;
		data_a[20973]<=8'd105;
		data_a[20974]<=8'd109;
		data_a[20975]<=8'd117;
		data_a[20976]<=8'd122;
		data_a[20977]<=8'd122;
		data_a[20978]<=8'd122;
		data_a[20979]<=8'd124;
		data_a[20980]<=8'd123;
		data_a[20981]<=8'd116;
		data_a[20982]<=8'd112;
		data_a[20983]<=8'd105;
		data_a[20984]<=8'd85;
		data_a[20985]<=8'd64;
		data_a[20986]<=8'd74;
		data_a[20987]<=8'd66;
		data_a[20988]<=8'd75;
		data_a[20989]<=8'd78;
		data_a[20990]<=8'd82;
		data_a[20991]<=8'd80;
		data_a[20992]<=8'd60;
		data_a[20993]<=8'd68;
		data_a[20994]<=8'd109;
		data_a[20995]<=8'd97;
		data_a[20996]<=8'd94;
		data_a[20997]<=8'd93;
		data_a[20998]<=8'd89;
		data_a[20999]<=8'd87;
		data_a[21000]<=8'd254;
		data_a[21001]<=8'd85;
		data_a[21002]<=8'd88;
		data_a[21003]<=8'd91;
		data_a[21004]<=8'd79;
		data_a[21005]<=8'd62;
		data_a[21006]<=8'd59;
		data_a[21007]<=8'd67;
		data_a[21008]<=8'd62;
		data_a[21009]<=8'd209;
		data_a[21010]<=8'd168;
		data_a[21011]<=8'd200;
		data_a[21012]<=8'd206;
		data_a[21013]<=8'd131;
		data_a[21014]<=8'd65;
		data_a[21015]<=8'd73;
		data_a[21016]<=8'd61;
		data_a[21017]<=8'd73;
		data_a[21018]<=8'd65;
		data_a[21019]<=8'd61;
		data_a[21020]<=8'd61;
		data_a[21021]<=8'd57;
		data_a[21022]<=8'd196;
		data_a[21023]<=8'd223;
		data_a[21024]<=8'd178;
		data_a[21025]<=8'd195;
		data_a[21026]<=8'd217;
		data_a[21027]<=8'd204;
		data_a[21028]<=8'd190;
		data_a[21029]<=8'd131;
		data_a[21030]<=8'd172;
		data_a[21031]<=8'd157;
		data_a[21032]<=8'd141;
		data_a[21033]<=8'd135;
		data_a[21034]<=8'd128;
		data_a[21035]<=8'd125;
		data_a[21036]<=8'd120;
		data_a[21037]<=8'd118;
		data_a[21038]<=8'd111;
		data_a[21039]<=8'd103;
		data_a[21040]<=8'd101;
		data_a[21041]<=8'd99;
		data_a[21042]<=8'd98;
		data_a[21043]<=8'd94;
		data_a[21044]<=8'd91;
		data_a[21045]<=8'd84;
		data_a[21046]<=8'd85;
		data_a[21047]<=8'd85;
		data_a[21048]<=8'd88;
		data_a[21049]<=8'd86;
		data_a[21050]<=8'd88;
		data_a[21051]<=8'd92;
		data_a[21052]<=8'd94;
		data_a[21053]<=8'd96;
		data_a[21054]<=8'd102;
		data_a[21055]<=8'd110;
		data_a[21056]<=8'd123;
		data_a[21057]<=8'd142;
		data_a[21058]<=8'd116;
		data_a[21059]<=8'd104;
		data_a[21060]<=8'd86;
		data_a[21061]<=8'd72;
		data_a[21062]<=8'd167;
		data_a[21063]<=8'd163;
		data_a[21064]<=8'd243;
		data_a[21065]<=8'd236;
		data_a[21066]<=8'd241;
		data_a[21067]<=8'd237;
		data_a[21068]<=8'd235;
		data_a[21069]<=8'd234;
		data_a[21070]<=8'd237;
		data_a[21071]<=8'd230;
		data_a[21072]<=8'd235;
		data_a[21073]<=8'd233;
		data_a[21074]<=8'd233;
		data_a[21075]<=8'd233;
		data_a[21076]<=8'd232;
		data_a[21077]<=8'd234;
		data_a[21078]<=8'd237;
		data_a[21079]<=8'd237;
		data_a[21080]<=8'd239;
		data_a[21081]<=8'd237;
		data_a[21082]<=8'd238;
		data_a[21083]<=8'd239;
		data_a[21084]<=8'd238;
		data_a[21085]<=8'd239;
		data_a[21086]<=8'd241;
		data_a[21087]<=8'd239;
		data_a[21088]<=8'd240;
		data_a[21089]<=8'd238;
		data_a[21090]<=8'd236;
		data_a[21091]<=8'd237;
		data_a[21092]<=8'd246;
		data_a[21093]<=8'd244;
		data_a[21094]<=8'd241;
		data_a[21095]<=8'd239;
		data_a[21096]<=8'd238;
		data_a[21097]<=8'd125;
		data_a[21098]<=8'd52;
		data_a[21099]<=8'd45;
		data_a[21100]<=8'd60;
		data_a[21101]<=8'd52;
		data_a[21102]<=8'd47;
		data_a[21103]<=8'd60;
		data_a[21104]<=8'd50;
		data_a[21105]<=8'd55;
		data_a[21106]<=8'd56;
		data_a[21107]<=8'd64;
		data_a[21108]<=8'd69;
		data_a[21109]<=8'd69;
		data_a[21110]<=8'd72;
		data_a[21111]<=8'd68;
		data_a[21112]<=8'd81;
		data_a[21113]<=8'd70;
		data_a[21114]<=8'd83;
		data_a[21115]<=8'd84;
		data_a[21116]<=8'd87;
		data_a[21117]<=8'd90;
		data_a[21118]<=8'd91;
		data_a[21119]<=8'd94;
		data_a[21120]<=8'd97;
		data_a[21121]<=8'd106;
		data_a[21122]<=8'd106;
		data_a[21123]<=8'd105;
		data_a[21124]<=8'd114;
		data_a[21125]<=8'd122;
		data_a[21126]<=8'd123;
		data_a[21127]<=8'd123;
		data_a[21128]<=8'd122;
		data_a[21129]<=8'd126;
		data_a[21130]<=8'd123;
		data_a[21131]<=8'd116;
		data_a[21132]<=8'd112;
		data_a[21133]<=8'd103;
		data_a[21134]<=8'd86;
		data_a[21135]<=8'd67;
		data_a[21136]<=8'd76;
		data_a[21137]<=8'd82;
		data_a[21138]<=8'd69;
		data_a[21139]<=8'd74;
		data_a[21140]<=8'd74;
		data_a[21141]<=8'd56;
		data_a[21142]<=8'd41;
		data_a[21143]<=8'd46;
		data_a[21144]<=8'd95;
		data_a[21145]<=8'd96;
		data_a[21146]<=8'd91;
		data_a[21147]<=8'd89;
		data_a[21148]<=8'd91;
		data_a[21149]<=8'd90;
		data_a[21150]<=8'd253;
		data_a[21151]<=8'd90;
		data_a[21152]<=8'd102;
		data_a[21153]<=8'd100;
		data_a[21154]<=8'd94;
		data_a[21155]<=8'd76;
		data_a[21156]<=8'd61;
		data_a[21157]<=8'd77;
		data_a[21158]<=8'd61;
		data_a[21159]<=8'd253;
		data_a[21160]<=8'd149;
		data_a[21161]<=8'd182;
		data_a[21162]<=8'd153;
		data_a[21163]<=8'd58;
		data_a[21164]<=8'd69;
		data_a[21165]<=8'd64;
		data_a[21166]<=8'd64;
		data_a[21167]<=8'd62;
		data_a[21168]<=8'd73;
		data_a[21169]<=8'd64;
		data_a[21170]<=8'd57;
		data_a[21171]<=8'd59;
		data_a[21172]<=8'd213;
		data_a[21173]<=8'd206;
		data_a[21174]<=8'd210;
		data_a[21175]<=8'd212;
		data_a[21176]<=8'd209;
		data_a[21177]<=8'd197;
		data_a[21178]<=8'd193;
		data_a[21179]<=8'd187;
		data_a[21180]<=8'd154;
		data_a[21181]<=8'd151;
		data_a[21182]<=8'd141;
		data_a[21183]<=8'd134;
		data_a[21184]<=8'd126;
		data_a[21185]<=8'd125;
		data_a[21186]<=8'd120;
		data_a[21187]<=8'd118;
		data_a[21188]<=8'd112;
		data_a[21189]<=8'd108;
		data_a[21190]<=8'd108;
		data_a[21191]<=8'd102;
		data_a[21192]<=8'd94;
		data_a[21193]<=8'd90;
		data_a[21194]<=8'd96;
		data_a[21195]<=8'd93;
		data_a[21196]<=8'd96;
		data_a[21197]<=8'd88;
		data_a[21198]<=8'd93;
		data_a[21199]<=8'd90;
		data_a[21200]<=8'd88;
		data_a[21201]<=8'd90;
		data_a[21202]<=8'd93;
		data_a[21203]<=8'd96;
		data_a[21204]<=8'd101;
		data_a[21205]<=8'd105;
		data_a[21206]<=8'd117;
		data_a[21207]<=8'd146;
		data_a[21208]<=8'd88;
		data_a[21209]<=8'd81;
		data_a[21210]<=8'd76;
		data_a[21211]<=8'd85;
		data_a[21212]<=8'd146;
		data_a[21213]<=8'd148;
		data_a[21214]<=8'd188;
		data_a[21215]<=8'd198;
		data_a[21216]<=8'd198;
		data_a[21217]<=8'd242;
		data_a[21218]<=8'd238;
		data_a[21219]<=8'd235;
		data_a[21220]<=8'd230;
		data_a[21221]<=8'd239;
		data_a[21222]<=8'd233;
		data_a[21223]<=8'd231;
		data_a[21224]<=8'd232;
		data_a[21225]<=8'd233;
		data_a[21226]<=8'd231;
		data_a[21227]<=8'd234;
		data_a[21228]<=8'd237;
		data_a[21229]<=8'd238;
		data_a[21230]<=8'd239;
		data_a[21231]<=8'd237;
		data_a[21232]<=8'd238;
		data_a[21233]<=8'd239;
		data_a[21234]<=8'd238;
		data_a[21235]<=8'd239;
		data_a[21236]<=8'd240;
		data_a[21237]<=8'd239;
		data_a[21238]<=8'd239;
		data_a[21239]<=8'd237;
		data_a[21240]<=8'd235;
		data_a[21241]<=8'd235;
		data_a[21242]<=8'd245;
		data_a[21243]<=8'd241;
		data_a[21244]<=8'd238;
		data_a[21245]<=8'd238;
		data_a[21246]<=8'd241;
		data_a[21247]<=8'd73;
		data_a[21248]<=8'd60;
		data_a[21249]<=8'd52;
		data_a[21250]<=8'd54;
		data_a[21251]<=8'd74;
		data_a[21252]<=8'd92;
		data_a[21253]<=8'd75;
		data_a[21254]<=8'd94;
		data_a[21255]<=8'd89;
		data_a[21256]<=8'd88;
		data_a[21257]<=8'd80;
		data_a[21258]<=8'd76;
		data_a[21259]<=8'd79;
		data_a[21260]<=8'd80;
		data_a[21261]<=8'd88;
		data_a[21262]<=8'd83;
		data_a[21263]<=8'd84;
		data_a[21264]<=8'd93;
		data_a[21265]<=8'd95;
		data_a[21266]<=8'd91;
		data_a[21267]<=8'd99;
		data_a[21268]<=8'd94;
		data_a[21269]<=8'd100;
		data_a[21270]<=8'd98;
		data_a[21271]<=8'd109;
		data_a[21272]<=8'd108;
		data_a[21273]<=8'd106;
		data_a[21274]<=8'd117;
		data_a[21275]<=8'd125;
		data_a[21276]<=8'd123;
		data_a[21277]<=8'd124;
		data_a[21278]<=8'd122;
		data_a[21279]<=8'd126;
		data_a[21280]<=8'd120;
		data_a[21281]<=8'd114;
		data_a[21282]<=8'd110;
		data_a[21283]<=8'd99;
		data_a[21284]<=8'd84;
		data_a[21285]<=8'd69;
		data_a[21286]<=8'd77;
		data_a[21287]<=8'd101;
		data_a[21288]<=8'd61;
		data_a[21289]<=8'd75;
		data_a[21290]<=8'd68;
		data_a[21291]<=8'd36;
		data_a[21292]<=8'd49;
		data_a[21293]<=8'd47;
		data_a[21294]<=8'd80;
		data_a[21295]<=8'd93;
		data_a[21296]<=8'd90;
		data_a[21297]<=8'd89;
		data_a[21298]<=8'd93;
		data_a[21299]<=8'd93;
		data_a[21300]<=8'd254;
		data_a[21301]<=8'd114;
		data_a[21302]<=8'd99;
		data_a[21303]<=8'd92;
		data_a[21304]<=8'd87;
		data_a[21305]<=8'd92;
		data_a[21306]<=8'd103;
		data_a[21307]<=8'd99;
		data_a[21308]<=8'd90;
		data_a[21309]<=8'd253;
		data_a[21310]<=8'd118;
		data_a[21311]<=8'd187;
		data_a[21312]<=8'd73;
		data_a[21313]<=8'd63;
		data_a[21314]<=8'd61;
		data_a[21315]<=8'd64;
		data_a[21316]<=8'd57;
		data_a[21317]<=8'd59;
		data_a[21318]<=8'd66;
		data_a[21319]<=8'd66;
		data_a[21320]<=8'd64;
		data_a[21321]<=8'd66;
		data_a[21322]<=8'd115;
		data_a[21323]<=8'd201;
		data_a[21324]<=8'd208;
		data_a[21325]<=8'd200;
		data_a[21326]<=8'd204;
		data_a[21327]<=8'd193;
		data_a[21328]<=8'd188;
		data_a[21329]<=8'd186;
		data_a[21330]<=8'd168;
		data_a[21331]<=8'd148;
		data_a[21332]<=8'd139;
		data_a[21333]<=8'd135;
		data_a[21334]<=8'd128;
		data_a[21335]<=8'd126;
		data_a[21336]<=8'd118;
		data_a[21337]<=8'd118;
		data_a[21338]<=8'd115;
		data_a[21339]<=8'd114;
		data_a[21340]<=8'd106;
		data_a[21341]<=8'd104;
		data_a[21342]<=8'd103;
		data_a[21343]<=8'd98;
		data_a[21344]<=8'd97;
		data_a[21345]<=8'd95;
		data_a[21346]<=8'd94;
		data_a[21347]<=8'd93;
		data_a[21348]<=8'd92;
		data_a[21349]<=8'd91;
		data_a[21350]<=8'd92;
		data_a[21351]<=8'd95;
		data_a[21352]<=8'd96;
		data_a[21353]<=8'd96;
		data_a[21354]<=8'd101;
		data_a[21355]<=8'd106;
		data_a[21356]<=8'd117;
		data_a[21357]<=8'd136;
		data_a[21358]<=8'd68;
		data_a[21359]<=8'd62;
		data_a[21360]<=8'd54;
		data_a[21361]<=8'd162;
		data_a[21362]<=8'd135;
		data_a[21363]<=8'd130;
		data_a[21364]<=8'd131;
		data_a[21365]<=8'd195;
		data_a[21366]<=8'd173;
		data_a[21367]<=8'd210;
		data_a[21368]<=8'd234;
		data_a[21369]<=8'd232;
		data_a[21370]<=8'd234;
		data_a[21371]<=8'd235;
		data_a[21372]<=8'd233;
		data_a[21373]<=8'd231;
		data_a[21374]<=8'd231;
		data_a[21375]<=8'd232;
		data_a[21376]<=8'd231;
		data_a[21377]<=8'd234;
		data_a[21378]<=8'd237;
		data_a[21379]<=8'd237;
		data_a[21380]<=8'd239;
		data_a[21381]<=8'd237;
		data_a[21382]<=8'd238;
		data_a[21383]<=8'd239;
		data_a[21384]<=8'd237;
		data_a[21385]<=8'd238;
		data_a[21386]<=8'd239;
		data_a[21387]<=8'd238;
		data_a[21388]<=8'd237;
		data_a[21389]<=8'd236;
		data_a[21390]<=8'd235;
		data_a[21391]<=8'd234;
		data_a[21392]<=8'd242;
		data_a[21393]<=8'd238;
		data_a[21394]<=8'd237;
		data_a[21395]<=8'd240;
		data_a[21396]<=8'd232;
		data_a[21397]<=8'd73;
		data_a[21398]<=8'd55;
		data_a[21399]<=8'd63;
		data_a[21400]<=8'd44;
		data_a[21401]<=8'd56;
		data_a[21402]<=8'd90;
		data_a[21403]<=8'd95;
		data_a[21404]<=8'd98;
		data_a[21405]<=8'd92;
		data_a[21406]<=8'd93;
		data_a[21407]<=8'd88;
		data_a[21408]<=8'd88;
		data_a[21409]<=8'd89;
		data_a[21410]<=8'd82;
		data_a[21411]<=8'd82;
		data_a[21412]<=8'd82;
		data_a[21413]<=8'd92;
		data_a[21414]<=8'd94;
		data_a[21415]<=8'd94;
		data_a[21416]<=8'd98;
		data_a[21417]<=8'd105;
		data_a[21418]<=8'd97;
		data_a[21419]<=8'd104;
		data_a[21420]<=8'd103;
		data_a[21421]<=8'd108;
		data_a[21422]<=8'd109;
		data_a[21423]<=8'd111;
		data_a[21424]<=8'd118;
		data_a[21425]<=8'd123;
		data_a[21426]<=8'd123;
		data_a[21427]<=8'd123;
		data_a[21428]<=8'd120;
		data_a[21429]<=8'd122;
		data_a[21430]<=8'd114;
		data_a[21431]<=8'd110;
		data_a[21432]<=8'd108;
		data_a[21433]<=8'd95;
		data_a[21434]<=8'd82;
		data_a[21435]<=8'd70;
		data_a[21436]<=8'd75;
		data_a[21437]<=8'd87;
		data_a[21438]<=8'd70;
		data_a[21439]<=8'd76;
		data_a[21440]<=8'd63;
		data_a[21441]<=8'd46;
		data_a[21442]<=8'd43;
		data_a[21443]<=8'd48;
		data_a[21444]<=8'd74;
		data_a[21445]<=8'd91;
		data_a[21446]<=8'd92;
		data_a[21447]<=8'd94;
		data_a[21448]<=8'd92;
		data_a[21449]<=8'd91;
		data_a[21450]<=8'd254;
		data_a[21451]<=8'd89;
		data_a[21452]<=8'd90;
		data_a[21453]<=8'd90;
		data_a[21454]<=8'd76;
		data_a[21455]<=8'd90;
		data_a[21456]<=8'd84;
		data_a[21457]<=8'd85;
		data_a[21458]<=8'd251;
		data_a[21459]<=8'd190;
		data_a[21460]<=8'd145;
		data_a[21461]<=8'd110;
		data_a[21462]<=8'd45;
		data_a[21463]<=8'd58;
		data_a[21464]<=8'd53;
		data_a[21465]<=8'd53;
		data_a[21466]<=8'd50;
		data_a[21467]<=8'd47;
		data_a[21468]<=8'd55;
		data_a[21469]<=8'd61;
		data_a[21470]<=8'd62;
		data_a[21471]<=8'd57;
		data_a[21472]<=8'd59;
		data_a[21473]<=8'd187;
		data_a[21474]<=8'd193;
		data_a[21475]<=8'd204;
		data_a[21476]<=8'd199;
		data_a[21477]<=8'd189;
		data_a[21478]<=8'd195;
		data_a[21479]<=8'd180;
		data_a[21480]<=8'd175;
		data_a[21481]<=8'd143;
		data_a[21482]<=8'd137;
		data_a[21483]<=8'd134;
		data_a[21484]<=8'd128;
		data_a[21485]<=8'd127;
		data_a[21486]<=8'd120;
		data_a[21487]<=8'd123;
		data_a[21488]<=8'd117;
		data_a[21489]<=8'd112;
		data_a[21490]<=8'd109;
		data_a[21491]<=8'd103;
		data_a[21492]<=8'd103;
		data_a[21493]<=8'd100;
		data_a[21494]<=8'd97;
		data_a[21495]<=8'd102;
		data_a[21496]<=8'd93;
		data_a[21497]<=8'd98;
		data_a[21498]<=8'd96;
		data_a[21499]<=8'd92;
		data_a[21500]<=8'd90;
		data_a[21501]<=8'd93;
		data_a[21502]<=8'd94;
		data_a[21503]<=8'd95;
		data_a[21504]<=8'd100;
		data_a[21505]<=8'd108;
		data_a[21506]<=8'd119;
		data_a[21507]<=8'd133;
		data_a[21508]<=8'd144;
		data_a[21509]<=8'd81;
		data_a[21510]<=8'd154;
		data_a[21511]<=8'd124;
		data_a[21512]<=8'd118;
		data_a[21513]<=8'd112;
		data_a[21514]<=8'd173;
		data_a[21515]<=8'd147;
		data_a[21516]<=8'd171;
		data_a[21517]<=8'd184;
		data_a[21518]<=8'd236;
		data_a[21519]<=8'd234;
		data_a[21520]<=8'd239;
		data_a[21521]<=8'd233;
		data_a[21522]<=8'd234;
		data_a[21523]<=8'd231;
		data_a[21524]<=8'd231;
		data_a[21525]<=8'd232;
		data_a[21526]<=8'd231;
		data_a[21527]<=8'd234;
		data_a[21528]<=8'd236;
		data_a[21529]<=8'd236;
		data_a[21530]<=8'd238;
		data_a[21531]<=8'd237;
		data_a[21532]<=8'd238;
		data_a[21533]<=8'd238;
		data_a[21534]<=8'd237;
		data_a[21535]<=8'd237;
		data_a[21536]<=8'd238;
		data_a[21537]<=8'd237;
		data_a[21538]<=8'd237;
		data_a[21539]<=8'd237;
		data_a[21540]<=8'd236;
		data_a[21541]<=8'd234;
		data_a[21542]<=8'd242;
		data_a[21543]<=8'd238;
		data_a[21544]<=8'd238;
		data_a[21545]<=8'd243;
		data_a[21546]<=8'd94;
		data_a[21547]<=8'd56;
		data_a[21548]<=8'd47;
		data_a[21549]<=8'd54;
		data_a[21550]<=8'd101;
		data_a[21551]<=8'd94;
		data_a[21552]<=8'd105;
		data_a[21553]<=8'd102;
		data_a[21554]<=8'd97;
		data_a[21555]<=8'd101;
		data_a[21556]<=8'd97;
		data_a[21557]<=8'd96;
		data_a[21558]<=8'd90;
		data_a[21559]<=8'd85;
		data_a[21560]<=8'd92;
		data_a[21561]<=8'd93;
		data_a[21562]<=8'd98;
		data_a[21563]<=8'd93;
		data_a[21564]<=8'd97;
		data_a[21565]<=8'd94;
		data_a[21566]<=8'd98;
		data_a[21567]<=8'd102;
		data_a[21568]<=8'd107;
		data_a[21569]<=8'd105;
		data_a[21570]<=8'd110;
		data_a[21571]<=8'd108;
		data_a[21572]<=8'd112;
		data_a[21573]<=8'd117;
		data_a[21574]<=8'd119;
		data_a[21575]<=8'd121;
		data_a[21576]<=8'd123;
		data_a[21577]<=8'd122;
		data_a[21578]<=8'd119;
		data_a[21579]<=8'd120;
		data_a[21580]<=8'd110;
		data_a[21581]<=8'd109;
		data_a[21582]<=8'd108;
		data_a[21583]<=8'd95;
		data_a[21584]<=8'd82;
		data_a[21585]<=8'd72;
		data_a[21586]<=8'd73;
		data_a[21587]<=8'd74;
		data_a[21588]<=8'd67;
		data_a[21589]<=8'd70;
		data_a[21590]<=8'd54;
		data_a[21591]<=8'd47;
		data_a[21592]<=8'd40;
		data_a[21593]<=8'd43;
		data_a[21594]<=8'd74;
		data_a[21595]<=8'd88;
		data_a[21596]<=8'd93;
		data_a[21597]<=8'd98;
		data_a[21598]<=8'd89;
		data_a[21599]<=8'd86;
		data_a[21600]<=8'd254;
		data_a[21601]<=8'd80;
		data_a[21602]<=8'd83;
		data_a[21603]<=8'd85;
		data_a[21604]<=8'd79;
		data_a[21605]<=8'd79;
		data_a[21606]<=8'd78;
		data_a[21607]<=8'd76;
		data_a[21608]<=8'd237;
		data_a[21609]<=8'd121;
		data_a[21610]<=8'd129;
		data_a[21611]<=8'd68;
		data_a[21612]<=8'd58;
		data_a[21613]<=8'd45;
		data_a[21614]<=8'd47;
		data_a[21615]<=8'd46;
		data_a[21616]<=8'd46;
		data_a[21617]<=8'd45;
		data_a[21618]<=8'd47;
		data_a[21619]<=8'd46;
		data_a[21620]<=8'd49;
		data_a[21621]<=8'd54;
		data_a[21622]<=8'd50;
		data_a[21623]<=8'd171;
		data_a[21624]<=8'd191;
		data_a[21625]<=8'd192;
		data_a[21626]<=8'd180;
		data_a[21627]<=8'd193;
		data_a[21628]<=8'd185;
		data_a[21629]<=8'd185;
		data_a[21630]<=8'd167;
		data_a[21631]<=8'd163;
		data_a[21632]<=8'd152;
		data_a[21633]<=8'd126;
		data_a[21634]<=8'd124;
		data_a[21635]<=8'd130;
		data_a[21636]<=8'd120;
		data_a[21637]<=8'd122;
		data_a[21638]<=8'd120;
		data_a[21639]<=8'd114;
		data_a[21640]<=8'd108;
		data_a[21641]<=8'd104;
		data_a[21642]<=8'd102;
		data_a[21643]<=8'd104;
		data_a[21644]<=8'd105;
		data_a[21645]<=8'd101;
		data_a[21646]<=8'd97;
		data_a[21647]<=8'd94;
		data_a[21648]<=8'd90;
		data_a[21649]<=8'd91;
		data_a[21650]<=8'd94;
		data_a[21651]<=8'd93;
		data_a[21652]<=8'd96;
		data_a[21653]<=8'd100;
		data_a[21654]<=8'd98;
		data_a[21655]<=8'd110;
		data_a[21656]<=8'd119;
		data_a[21657]<=8'd132;
		data_a[21658]<=8'd148;
		data_a[21659]<=8'd91;
		data_a[21660]<=8'd117;
		data_a[21661]<=8'd108;
		data_a[21662]<=8'd107;
		data_a[21663]<=8'd120;
		data_a[21664]<=8'd144;
		data_a[21665]<=8'd160;
		data_a[21666]<=8'd182;
		data_a[21667]<=8'd195;
		data_a[21668]<=8'd203;
		data_a[21669]<=8'd219;
		data_a[21670]<=8'd242;
		data_a[21671]<=8'd230;
		data_a[21672]<=8'd230;
		data_a[21673]<=8'd234;
		data_a[21674]<=8'd228;
		data_a[21675]<=8'd227;
		data_a[21676]<=8'd230;
		data_a[21677]<=8'd237;
		data_a[21678]<=8'd237;
		data_a[21679]<=8'd235;
		data_a[21680]<=8'd238;
		data_a[21681]<=8'd239;
		data_a[21682]<=8'd237;
		data_a[21683]<=8'd239;
		data_a[21684]<=8'd238;
		data_a[21685]<=8'd237;
		data_a[21686]<=8'd239;
		data_a[21687]<=8'd238;
		data_a[21688]<=8'd238;
		data_a[21689]<=8'd236;
		data_a[21690]<=8'd230;
		data_a[21691]<=8'd236;
		data_a[21692]<=8'd242;
		data_a[21693]<=8'd238;
		data_a[21694]<=8'd238;
		data_a[21695]<=8'd239;
		data_a[21696]<=8'd71;
		data_a[21697]<=8'd59;
		data_a[21698]<=8'd46;
		data_a[21699]<=8'd49;
		data_a[21700]<=8'd88;
		data_a[21701]<=8'd102;
		data_a[21702]<=8'd106;
		data_a[21703]<=8'd103;
		data_a[21704]<=8'd102;
		data_a[21705]<=8'd100;
		data_a[21706]<=8'd101;
		data_a[21707]<=8'd98;
		data_a[21708]<=8'd95;
		data_a[21709]<=8'd94;
		data_a[21710]<=8'd92;
		data_a[21711]<=8'd93;
		data_a[21712]<=8'd95;
		data_a[21713]<=8'd96;
		data_a[21714]<=8'd100;
		data_a[21715]<=8'd104;
		data_a[21716]<=8'd107;
		data_a[21717]<=8'd108;
		data_a[21718]<=8'd109;
		data_a[21719]<=8'd110;
		data_a[21720]<=8'd113;
		data_a[21721]<=8'd114;
		data_a[21722]<=8'd115;
		data_a[21723]<=8'd118;
		data_a[21724]<=8'd122;
		data_a[21725]<=8'd124;
		data_a[21726]<=8'd124;
		data_a[21727]<=8'd121;
		data_a[21728]<=8'd118;
		data_a[21729]<=8'd115;
		data_a[21730]<=8'd109;
		data_a[21731]<=8'd109;
		data_a[21732]<=8'd103;
		data_a[21733]<=8'd90;
		data_a[21734]<=8'd82;
		data_a[21735]<=8'd70;
		data_a[21736]<=8'd72;
		data_a[21737]<=8'd80;
		data_a[21738]<=8'd70;
		data_a[21739]<=8'd66;
		data_a[21740]<=8'd44;
		data_a[21741]<=8'd46;
		data_a[21742]<=8'd53;
		data_a[21743]<=8'd48;
		data_a[21744]<=8'd81;
		data_a[21745]<=8'd88;
		data_a[21746]<=8'd94;
		data_a[21747]<=8'd93;
		data_a[21748]<=8'd90;
		data_a[21749]<=8'd88;
		data_a[21750]<=8'd254;
		data_a[21751]<=8'd79;
		data_a[21752]<=8'd73;
		data_a[21753]<=8'd80;
		data_a[21754]<=8'd77;
		data_a[21755]<=8'd76;
		data_a[21756]<=8'd74;
		data_a[21757]<=8'd147;
		data_a[21758]<=8'd253;
		data_a[21759]<=8'd130;
		data_a[21760]<=8'd69;
		data_a[21761]<=8'd55;
		data_a[21762]<=8'd75;
		data_a[21763]<=8'd39;
		data_a[21764]<=8'd37;
		data_a[21765]<=8'd41;
		data_a[21766]<=8'd39;
		data_a[21767]<=8'd39;
		data_a[21768]<=8'd42;
		data_a[21769]<=8'd40;
		data_a[21770]<=8'd44;
		data_a[21771]<=8'd51;
		data_a[21772]<=8'd52;
		data_a[21773]<=8'd154;
		data_a[21774]<=8'd184;
		data_a[21775]<=8'd191;
		data_a[21776]<=8'd192;
		data_a[21777]<=8'd186;
		data_a[21778]<=8'd189;
		data_a[21779]<=8'd180;
		data_a[21780]<=8'd169;
		data_a[21781]<=8'd147;
		data_a[21782]<=8'd149;
		data_a[21783]<=8'd153;
		data_a[21784]<=8'd142;
		data_a[21785]<=8'd117;
		data_a[21786]<=8'd113;
		data_a[21787]<=8'd125;
		data_a[21788]<=8'd120;
		data_a[21789]<=8'd113;
		data_a[21790]<=8'd106;
		data_a[21791]<=8'd103;
		data_a[21792]<=8'd101;
		data_a[21793]<=8'd103;
		data_a[21794]<=8'd104;
		data_a[21795]<=8'd102;
		data_a[21796]<=8'd99;
		data_a[21797]<=8'd98;
		data_a[21798]<=8'd93;
		data_a[21799]<=8'd97;
		data_a[21800]<=8'd94;
		data_a[21801]<=8'd99;
		data_a[21802]<=8'd101;
		data_a[21803]<=8'd96;
		data_a[21804]<=8'd101;
		data_a[21805]<=8'd109;
		data_a[21806]<=8'd118;
		data_a[21807]<=8'd127;
		data_a[21808]<=8'd139;
		data_a[21809]<=8'd110;
		data_a[21810]<=8'd107;
		data_a[21811]<=8'd102;
		data_a[21812]<=8'd106;
		data_a[21813]<=8'd148;
		data_a[21814]<=8'd142;
		data_a[21815]<=8'd179;
		data_a[21816]<=8'd178;
		data_a[21817]<=8'd178;
		data_a[21818]<=8'd170;
		data_a[21819]<=8'd175;
		data_a[21820]<=8'd179;
		data_a[21821]<=8'd235;
		data_a[21822]<=8'd234;
		data_a[21823]<=8'd230;
		data_a[21824]<=8'd230;
		data_a[21825]<=8'd231;
		data_a[21826]<=8'd231;
		data_a[21827]<=8'd233;
		data_a[21828]<=8'd234;
		data_a[21829]<=8'd237;
		data_a[21830]<=8'd232;
		data_a[21831]<=8'd239;
		data_a[21832]<=8'd245;
		data_a[21833]<=8'd242;
		data_a[21834]<=8'd246;
		data_a[21835]<=8'd235;
		data_a[21836]<=8'd233;
		data_a[21837]<=8'd241;
		data_a[21838]<=8'd235;
		data_a[21839]<=8'd240;
		data_a[21840]<=8'd237;
		data_a[21841]<=8'd231;
		data_a[21842]<=8'd237;
		data_a[21843]<=8'd242;
		data_a[21844]<=8'd240;
		data_a[21845]<=8'd165;
		data_a[21846]<=8'd76;
		data_a[21847]<=8'd60;
		data_a[21848]<=8'd51;
		data_a[21849]<=8'd43;
		data_a[21850]<=8'd88;
		data_a[21851]<=8'd98;
		data_a[21852]<=8'd107;
		data_a[21853]<=8'd108;
		data_a[21854]<=8'd104;
		data_a[21855]<=8'd103;
		data_a[21856]<=8'd104;
		data_a[21857]<=8'd101;
		data_a[21858]<=8'd98;
		data_a[21859]<=8'd97;
		data_a[21860]<=8'd94;
		data_a[21861]<=8'd96;
		data_a[21862]<=8'd100;
		data_a[21863]<=8'd99;
		data_a[21864]<=8'd101;
		data_a[21865]<=8'd105;
		data_a[21866]<=8'd109;
		data_a[21867]<=8'd111;
		data_a[21868]<=8'd112;
		data_a[21869]<=8'd112;
		data_a[21870]<=8'd113;
		data_a[21871]<=8'd114;
		data_a[21872]<=8'd115;
		data_a[21873]<=8'd117;
		data_a[21874]<=8'd120;
		data_a[21875]<=8'd122;
		data_a[21876]<=8'd121;
		data_a[21877]<=8'd119;
		data_a[21878]<=8'd118;
		data_a[21879]<=8'd115;
		data_a[21880]<=8'd109;
		data_a[21881]<=8'd107;
		data_a[21882]<=8'd101;
		data_a[21883]<=8'd91;
		data_a[21884]<=8'd84;
		data_a[21885]<=8'd72;
		data_a[21886]<=8'd71;
		data_a[21887]<=8'd87;
		data_a[21888]<=8'd107;
		data_a[21889]<=8'd59;
		data_a[21890]<=8'd39;
		data_a[21891]<=8'd48;
		data_a[21892]<=8'd57;
		data_a[21893]<=8'd52;
		data_a[21894]<=8'd85;
		data_a[21895]<=8'd89;
		data_a[21896]<=8'd93;
		data_a[21897]<=8'd93;
		data_a[21898]<=8'd91;
		data_a[21899]<=8'd89;
		data_a[21900]<=8'd254;
		data_a[21901]<=8'd76;
		data_a[21902]<=8'd79;
		data_a[21903]<=8'd74;
		data_a[21904]<=8'd87;
		data_a[21905]<=8'd89;
		data_a[21906]<=8'd59;
		data_a[21907]<=8'd243;
		data_a[21908]<=8'd215;
		data_a[21909]<=8'd94;
		data_a[21910]<=8'd68;
		data_a[21911]<=8'd67;
		data_a[21912]<=8'd63;
		data_a[21913]<=8'd37;
		data_a[21914]<=8'd59;
		data_a[21915]<=8'd43;
		data_a[21916]<=8'd54;
		data_a[21917]<=8'd52;
		data_a[21918]<=8'd53;
		data_a[21919]<=8'd45;
		data_a[21920]<=8'd42;
		data_a[21921]<=8'd43;
		data_a[21922]<=8'd43;
		data_a[21923]<=8'd109;
		data_a[21924]<=8'd166;
		data_a[21925]<=8'd179;
		data_a[21926]<=8'd184;
		data_a[21927]<=8'd181;
		data_a[21928]<=8'd199;
		data_a[21929]<=8'd171;
		data_a[21930]<=8'd162;
		data_a[21931]<=8'd157;
		data_a[21932]<=8'd146;
		data_a[21933]<=8'd144;
		data_a[21934]<=8'd142;
		data_a[21935]<=8'd141;
		data_a[21936]<=8'd140;
		data_a[21937]<=8'd120;
		data_a[21938]<=8'd107;
		data_a[21939]<=8'd118;
		data_a[21940]<=8'd111;
		data_a[21941]<=8'd107;
		data_a[21942]<=8'd104;
		data_a[21943]<=8'd103;
		data_a[21944]<=8'd102;
		data_a[21945]<=8'd99;
		data_a[21946]<=8'd96;
		data_a[21947]<=8'd95;
		data_a[21948]<=8'd95;
		data_a[21949]<=8'd94;
		data_a[21950]<=8'd92;
		data_a[21951]<=8'd93;
		data_a[21952]<=8'd95;
		data_a[21953]<=8'd94;
		data_a[21954]<=8'd102;
		data_a[21955]<=8'd113;
		data_a[21956]<=8'd117;
		data_a[21957]<=8'd129;
		data_a[21958]<=8'd118;
		data_a[21959]<=8'd104;
		data_a[21960]<=8'd92;
		data_a[21961]<=8'd85;
		data_a[21962]<=8'd126;
		data_a[21963]<=8'd129;
		data_a[21964]<=8'd151;
		data_a[21965]<=8'd140;
		data_a[21966]<=8'd138;
		data_a[21967]<=8'd144;
		data_a[21968]<=8'd146;
		data_a[21969]<=8'd151;
		data_a[21970]<=8'd161;
		data_a[21971]<=8'd239;
		data_a[21972]<=8'd232;
		data_a[21973]<=8'd231;
		data_a[21974]<=8'd223;
		data_a[21975]<=8'd233;
		data_a[21976]<=8'd238;
		data_a[21977]<=8'd224;
		data_a[21978]<=8'd237;
		data_a[21979]<=8'd233;
		data_a[21980]<=8'd240;
		data_a[21981]<=8'd232;
		data_a[21982]<=8'd229;
		data_a[21983]<=8'd233;
		data_a[21984]<=8'd219;
		data_a[21985]<=8'd241;
		data_a[21986]<=8'd236;
		data_a[21987]<=8'd237;
		data_a[21988]<=8'd233;
		data_a[21989]<=8'd233;
		data_a[21990]<=8'd236;
		data_a[21991]<=8'd232;
		data_a[21992]<=8'd238;
		data_a[21993]<=8'd242;
		data_a[21994]<=8'd243;
		data_a[21995]<=8'd100;
		data_a[21996]<=8'd72;
		data_a[21997]<=8'd57;
		data_a[21998]<=8'd52;
		data_a[21999]<=8'd44;
		data_a[22000]<=8'd80;
		data_a[22001]<=8'd99;
		data_a[22002]<=8'd106;
		data_a[22003]<=8'd109;
		data_a[22004]<=8'd106;
		data_a[22005]<=8'd105;
		data_a[22006]<=8'd106;
		data_a[22007]<=8'd103;
		data_a[22008]<=8'd101;
		data_a[22009]<=8'd100;
		data_a[22010]<=8'd97;
		data_a[22011]<=8'd98;
		data_a[22012]<=8'd101;
		data_a[22013]<=8'd101;
		data_a[22014]<=8'd103;
		data_a[22015]<=8'd107;
		data_a[22016]<=8'd111;
		data_a[22017]<=8'd113;
		data_a[22018]<=8'd112;
		data_a[22019]<=8'd112;
		data_a[22020]<=8'd114;
		data_a[22021]<=8'd115;
		data_a[22022]<=8'd117;
		data_a[22023]<=8'd118;
		data_a[22024]<=8'd120;
		data_a[22025]<=8'd121;
		data_a[22026]<=8'd120;
		data_a[22027]<=8'd119;
		data_a[22028]<=8'd117;
		data_a[22029]<=8'd115;
		data_a[22030]<=8'd109;
		data_a[22031]<=8'd105;
		data_a[22032]<=8'd98;
		data_a[22033]<=8'd92;
		data_a[22034]<=8'd85;
		data_a[22035]<=8'd75;
		data_a[22036]<=8'd75;
		data_a[22037]<=8'd85;
		data_a[22038]<=8'd96;
		data_a[22039]<=8'd67;
		data_a[22040]<=8'd44;
		data_a[22041]<=8'd47;
		data_a[22042]<=8'd58;
		data_a[22043]<=8'd50;
		data_a[22044]<=8'd87;
		data_a[22045]<=8'd88;
		data_a[22046]<=8'd90;
		data_a[22047]<=8'd91;
		data_a[22048]<=8'd90;
		data_a[22049]<=8'd88;
		data_a[22050]<=8'd254;
		data_a[22051]<=8'd74;
		data_a[22052]<=8'd72;
		data_a[22053]<=8'd79;
		data_a[22054]<=8'd76;
		data_a[22055]<=8'd80;
		data_a[22056]<=8'd112;
		data_a[22057]<=8'd254;
		data_a[22058]<=8'd120;
		data_a[22059]<=8'd69;
		data_a[22060]<=8'd70;
		data_a[22061]<=8'd47;
		data_a[22062]<=8'd57;
		data_a[22063]<=8'd45;
		data_a[22064]<=8'd45;
		data_a[22065]<=8'd43;
		data_a[22066]<=8'd43;
		data_a[22067]<=8'd44;
		data_a[22068]<=8'd50;
		data_a[22069]<=8'd47;
		data_a[22070]<=8'd50;
		data_a[22071]<=8'd54;
		data_a[22072]<=8'd58;
		data_a[22073]<=8'd89;
		data_a[22074]<=8'd171;
		data_a[22075]<=8'd169;
		data_a[22076]<=8'd178;
		data_a[22077]<=8'd191;
		data_a[22078]<=8'd181;
		data_a[22079]<=8'd179;
		data_a[22080]<=8'd184;
		data_a[22081]<=8'd154;
		data_a[22082]<=8'd157;
		data_a[22083]<=8'd149;
		data_a[22084]<=8'd147;
		data_a[22085]<=8'd141;
		data_a[22086]<=8'd136;
		data_a[22087]<=8'd132;
		data_a[22088]<=8'd132;
		data_a[22089]<=8'd129;
		data_a[22090]<=8'd109;
		data_a[22091]<=8'd104;
		data_a[22092]<=8'd100;
		data_a[22093]<=8'd98;
		data_a[22094]<=8'd95;
		data_a[22095]<=8'd91;
		data_a[22096]<=8'd89;
		data_a[22097]<=8'd89;
		data_a[22098]<=8'd97;
		data_a[22099]<=8'd89;
		data_a[22100]<=8'd96;
		data_a[22101]<=8'd89;
		data_a[22102]<=8'd94;
		data_a[22103]<=8'd103;
		data_a[22104]<=8'd104;
		data_a[22105]<=8'd117;
		data_a[22106]<=8'd133;
		data_a[22107]<=8'd110;
		data_a[22108]<=8'd87;
		data_a[22109]<=8'd66;
		data_a[22110]<=8'd77;
		data_a[22111]<=8'd79;
		data_a[22112]<=8'd48;
		data_a[22113]<=8'd61;
		data_a[22114]<=8'd50;
		data_a[22115]<=8'd92;
		data_a[22116]<=8'd113;
		data_a[22117]<=8'd113;
		data_a[22118]<=8'd117;
		data_a[22119]<=8'd134;
		data_a[22120]<=8'd130;
		data_a[22121]<=8'd209;
		data_a[22122]<=8'd234;
		data_a[22123]<=8'd231;
		data_a[22124]<=8'd227;
		data_a[22125]<=8'd119;
		data_a[22126]<=8'd102;
		data_a[22127]<=8'd206;
		data_a[22128]<=8'd232;
		data_a[22129]<=8'd236;
		data_a[22130]<=8'd236;
		data_a[22131]<=8'd239;
		data_a[22132]<=8'd229;
		data_a[22133]<=8'd178;
		data_a[22134]<=8'd196;
		data_a[22135]<=8'd231;
		data_a[22136]<=8'd238;
		data_a[22137]<=8'd234;
		data_a[22138]<=8'd240;
		data_a[22139]<=8'd233;
		data_a[22140]<=8'd237;
		data_a[22141]<=8'd235;
		data_a[22142]<=8'd239;
		data_a[22143]<=8'd236;
		data_a[22144]<=8'd239;
		data_a[22145]<=8'd75;
		data_a[22146]<=8'd67;
		data_a[22147]<=8'd55;
		data_a[22148]<=8'd49;
		data_a[22149]<=8'd48;
		data_a[22150]<=8'd57;
		data_a[22151]<=8'd99;
		data_a[22152]<=8'd102;
		data_a[22153]<=8'd107;
		data_a[22154]<=8'd107;
		data_a[22155]<=8'd106;
		data_a[22156]<=8'd108;
		data_a[22157]<=8'd106;
		data_a[22158]<=8'd104;
		data_a[22159]<=8'd103;
		data_a[22160]<=8'd101;
		data_a[22161]<=8'd102;
		data_a[22162]<=8'd101;
		data_a[22163]<=8'd102;
		data_a[22164]<=8'd106;
		data_a[22165]<=8'd111;
		data_a[22166]<=8'd114;
		data_a[22167]<=8'd114;
		data_a[22168]<=8'd112;
		data_a[22169]<=8'd111;
		data_a[22170]<=8'd113;
		data_a[22171]<=8'd115;
		data_a[22172]<=8'd117;
		data_a[22173]<=8'd118;
		data_a[22174]<=8'd119;
		data_a[22175]<=8'd120;
		data_a[22176]<=8'd120;
		data_a[22177]<=8'd120;
		data_a[22178]<=8'd116;
		data_a[22179]<=8'd114;
		data_a[22180]<=8'd109;
		data_a[22181]<=8'd103;
		data_a[22182]<=8'd97;
		data_a[22183]<=8'd93;
		data_a[22184]<=8'd86;
		data_a[22185]<=8'd76;
		data_a[22186]<=8'd71;
		data_a[22187]<=8'd86;
		data_a[22188]<=8'd88;
		data_a[22189]<=8'd115;
		data_a[22190]<=8'd36;
		data_a[22191]<=8'd52;
		data_a[22192]<=8'd53;
		data_a[22193]<=8'd79;
		data_a[22194]<=8'd85;
		data_a[22195]<=8'd85;
		data_a[22196]<=8'd87;
		data_a[22197]<=8'd89;
		data_a[22198]<=8'd88;
		data_a[22199]<=8'd86;
		data_a[22200]<=8'd254;
		data_a[22201]<=8'd69;
		data_a[22202]<=8'd74;
		data_a[22203]<=8'd73;
		data_a[22204]<=8'd77;
		data_a[22205]<=8'd69;
		data_a[22206]<=8'd253;
		data_a[22207]<=8'd232;
		data_a[22208]<=8'd73;
		data_a[22209]<=8'd65;
		data_a[22210]<=8'd58;
		data_a[22211]<=8'd50;
		data_a[22212]<=8'd51;
		data_a[22213]<=8'd43;
		data_a[22214]<=8'd37;
		data_a[22215]<=8'd39;
		data_a[22216]<=8'd36;
		data_a[22217]<=8'd38;
		data_a[22218]<=8'd43;
		data_a[22219]<=8'd40;
		data_a[22220]<=8'd44;
		data_a[22221]<=8'd47;
		data_a[22222]<=8'd51;
		data_a[22223]<=8'd55;
		data_a[22224]<=8'd124;
		data_a[22225]<=8'd170;
		data_a[22226]<=8'd159;
		data_a[22227]<=8'd167;
		data_a[22228]<=8'd166;
		data_a[22229]<=8'd162;
		data_a[22230]<=8'd159;
		data_a[22231]<=8'd176;
		data_a[22232]<=8'd161;
		data_a[22233]<=8'd148;
		data_a[22234]<=8'd144;
		data_a[22235]<=8'd144;
		data_a[22236]<=8'd135;
		data_a[22237]<=8'd130;
		data_a[22238]<=8'd132;
		data_a[22239]<=8'd127;
		data_a[22240]<=8'd121;
		data_a[22241]<=8'd117;
		data_a[22242]<=8'd114;
		data_a[22243]<=8'd113;
		data_a[22244]<=8'd112;
		data_a[22245]<=8'd109;
		data_a[22246]<=8'd109;
		data_a[22247]<=8'd110;
		data_a[22248]<=8'd117;
		data_a[22249]<=8'd114;
		data_a[22250]<=8'd126;
		data_a[22251]<=8'd120;
		data_a[22252]<=8'd126;
		data_a[22253]<=8'd133;
		data_a[22254]<=8'd128;
		data_a[22255]<=8'd127;
		data_a[22256]<=8'd107;
		data_a[22257]<=8'd47;
		data_a[22258]<=8'd47;
		data_a[22259]<=8'd44;
		data_a[22260]<=8'd44;
		data_a[22261]<=8'd42;
		data_a[22262]<=8'd59;
		data_a[22263]<=8'd44;
		data_a[22264]<=8'd44;
		data_a[22265]<=8'd52;
		data_a[22266]<=8'd60;

	end
	
	// This block is activated at the positive edge of the writing clock (25MHz)
	// This block is responsible to write the datat in buffer port A
	always @(posedge w_clk) 
	begin
		// Check if the writing enable is activated or not to write on port B
		if(w_en_a)
		begin
			err_w_a <= 0;
			data_a[w_addr_a] <= d_in_a;
		end
		else
			err_w_a <= 1;
				
	end
	
	// This block is activated at the positive edge of the reading clock (50MHz)
	// This block is responsible to read from the port A and read and write from port B
	// Port B is read and writen at the same clock (50MHz) as it is read by VGA and writen by Sobel operator
	always @(posedge r_clk)
	begin
		d_out_a <= data_a[r_addr_a];		// Set the A out data from the registers of A
		d_out_b <= data_b[r_addr_b];		// Set the B out data from the registers of B
		
		// Check if the writing enable is activated or not to write on port B
		if(w_en_b == 1)
		begin
			err_w_b <= 0;
			data_b[w_addr_b] <= d_in_b;	// Store the input data
		end
		else
			err_w_b <= 1;
	end
	
endmodule
